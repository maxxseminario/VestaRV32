/home/mseminario2/chips/myshkin/ic/abstracts/myshkin_abs/GlitchFilter/GlitchFilter.lef