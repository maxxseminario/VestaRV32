/home/mseminario2/chips/myshkin/ic/abstracts/myshkin_abs/PowerOnResetCheng/PowerOnResetCheng.lef