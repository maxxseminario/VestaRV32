##
## LEF for PtnCells ;
## created by Innovus v20.12-s088_1 on Sat Nov  1 22:39:00 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MCU
  CLASS BLOCK ;
  SIZE 1186.000000 BY 686.000000 ;
  FOREIGN MCU 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN resetn_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.542 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 25.922 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 114.101 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6  ;
    ANTENNAMAXAREACAR 974.013 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 4292.32 LAYER M6  ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 131.365000 0.000000 131.465000 0.520000 ;
    END
  END resetn_in
  PIN resetn_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.325 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.474 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 111.130000 0.000000 111.230000 0.520000 ;
    END
  END resetn_out
  PIN resetn_dir
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.3585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6654 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 121.725000 0.000000 121.825000 0.520000 ;
    END
  END resetn_dir
  PIN resetn_ren
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.6965 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1086 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 125.685000 0.000000 125.785000 0.520000 ;
    END
  END resetn_ren
  PIN prt1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.495 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 583.026 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 2565.02 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 45.565000 1186.000000 45.665000 ;
    END
  END prt1_in[7]
  PIN prt1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1925 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.447 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 5.658 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9392 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 235.808 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1018.15 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 133.565000 1186.000000 133.665000 ;
    END
  END prt1_in[6]
  PIN prt1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0325 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.943 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 3.526 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5584 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3  ;
    ANTENNAMAXAREACAR 173.829 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 748.569 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 221.565000 1186.000000 221.665000 ;
    END
  END prt1_in[5]
  PIN prt1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.855 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 13.684 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.2976 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2577 LAYER M3  ;
    ANTENNAMAXAREACAR 64.8822 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 284.876 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.935444 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 309.565000 1186.000000 309.665000 ;
    END
  END prt1_in[4]
  PIN prt1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.176 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1936 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.52 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.848 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.964 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2364 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 19.36 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 21.648 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER M5  ;
    ANTENNAMAXAREACAR 146.799 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 177.903 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.88679 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 397.565000 1186.000000 397.665000 ;
    END
  END prt1_in[3]
  PIN prt1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0155 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.0682 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 11.178 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.2272 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 1.916 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5184 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1776 LAYER M4  ;
    ANTENNAMAXAREACAR 63.2544 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 281.931 LAYER M4  ;
    ANTENNAMAXCUTCAR 2.43902 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 485.565000 1186.000000 485.665000 ;
    END
  END prt1_in[2]
  PIN prt1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2935 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7354 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 3.092 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6928 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3  ;
    ANTENNAMAXAREACAR 37.9202 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 166.811 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 573.565000 1186.000000 573.665000 ;
    END
  END prt1_in[1]
  PIN prt1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8195 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.4058 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 4.662 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.5568 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3  ;
    ANTENNAMAXAREACAR 218.144 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 959.649 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 661.565000 1186.000000 661.665000 ;
    END
  END prt1_in[0]
  PIN prt1_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 8.214 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.1856 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 25.330000 1186.000000 25.430000 ;
    END
  END prt1_out[7]
  PIN prt1_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 113.330000 1186.000000 113.430000 ;
    END
  END prt1_out[6]
  PIN prt1_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 6.043 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.6772 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 201.330000 1186.000000 201.430000 ;
    END
  END prt1_out[5]
  PIN prt1_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 289.330000 1186.000000 289.430000 ;
    END
  END prt1_out[4]
  PIN prt1_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.976 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2944 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 8.742 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.5088 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 377.330000 1186.000000 377.430000 ;
    END
  END prt1_out[3]
  PIN prt1_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 465.330000 1186.000000 465.430000 ;
    END
  END prt1_out[2]
  PIN prt1_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 553.330000 1186.000000 553.430000 ;
    END
  END prt1_out[1]
  PIN prt1_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 10.699 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.1636 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 641.330000 1186.000000 641.430000 ;
    END
  END prt1_out[0]
  PIN prt1_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 35.925000 1186.000000 36.025000 ;
    END
  END prt1_dir[7]
  PIN prt1_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 123.925000 1186.000000 124.025000 ;
    END
  END prt1_dir[6]
  PIN prt1_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2345 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0758 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 9.306 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.9904 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 211.925000 1186.000000 212.025000 ;
    END
  END prt1_dir[5]
  PIN prt1_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 299.925000 1186.000000 300.025000 ;
    END
  END prt1_dir[4]
  PIN prt1_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7365 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2406 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 7.006 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8704 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 387.925000 1186.000000 388.025000 ;
    END
  END prt1_dir[3]
  PIN prt1_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2155 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9482 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 8.898 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.1952 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 475.925000 1186.000000 476.025000 ;
    END
  END prt1_dir[2]
  PIN prt1_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3486 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 563.925000 1186.000000 564.025000 ;
    END
  END prt1_dir[1]
  PIN prt1_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 11.5345 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.8398 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 651.925000 1186.000000 652.025000 ;
    END
  END prt1_dir[0]
  PIN prt1_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2262 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.426 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3184 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 39.885000 1186.000000 39.985000 ;
    END
  END prt1_ren[7]
  PIN prt1_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 13.4255 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.2042 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 127.885000 1186.000000 127.985000 ;
    END
  END prt1_ren[6]
  PIN prt1_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 215.885000 1186.000000 215.985000 ;
    END
  END prt1_ren[5]
  PIN prt1_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 303.885000 1186.000000 303.985000 ;
    END
  END prt1_ren[4]
  PIN prt1_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5302 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.802 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1728 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 391.885000 1186.000000 391.985000 ;
    END
  END prt1_ren[3]
  PIN prt1_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5655 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1322 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.522 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5408 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 479.885000 1186.000000 479.985000 ;
    END
  END prt1_ren[2]
  PIN prt1_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 11.5305 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.8222 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 567.885000 1186.000000 567.985000 ;
    END
  END prt1_ren[1]
  PIN prt1_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 11.5305 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.8222 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1185.480000 655.885000 1186.000000 655.985000 ;
    END
  END prt1_ren[0]
  PIN prt2_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7505 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3462 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0671 LAYER M2  ;
    ANTENNAMAXAREACAR 15.8756 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 68.1639 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.298063 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 302.965000 0.000000 303.065000 0.520000 ;
    END
  END prt2_in[7]
  PIN prt2_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5322 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2  ;
    ANTENNAMAXAREACAR 18.9193 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 83.7118 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 388.765000 0.000000 388.865000 0.520000 ;
    END
  END prt2_in[6]
  PIN prt2_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.731 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 2.282 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0848 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M3  ;
    ANTENNAMAXAREACAR 130.435 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 562.465 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.63265 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 474.565000 0.000000 474.665000 0.520000 ;
    END
  END prt2_in[5]
  PIN prt2_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7595 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3418 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 4.898 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5952 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3  ;
    ANTENNAMAXAREACAR 148.225 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 642.715 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 560.365000 0.000000 560.465000 0.520000 ;
    END
  END prt2_in[4]
  PIN prt2_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3916 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 2.64 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.08 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3816 LAYER M4  ;
    ANTENNAMAXAREACAR 8.48218 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 11.9754 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 646.165000 0.000000 646.265000 0.520000 ;
    END
  END prt2_in[3]
  PIN prt2_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 30.182 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 132.845 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3  ;
    ANTENNAMAXAREACAR 903.833 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 3969.24 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 731.965000 0.000000 732.065000 0.520000 ;
    END
  END prt2_in[2]
  PIN prt2_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.931 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0964 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 20.862 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.8368 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0451 LAYER M3  ;
    ANTENNAMAXAREACAR 479.446 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 2108.48 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.886918 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 817.765000 0.000000 817.865000 0.520000 ;
    END
  END prt2_in[1]
  PIN prt2_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5575 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.497 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M2  ;
    ANTENNAMAXAREACAR 3.38679 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 14.6436 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.104822 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 903.565000 0.000000 903.665000 0.520000 ;
    END
  END prt2_in[0]
  PIN prt2_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.471 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0724 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 9.582 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.2048 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 282.730000 0.000000 282.830000 0.520000 ;
    END
  END prt2_out[7]
  PIN prt2_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.721 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 368.530000 0.000000 368.630000 0.520000 ;
    END
  END prt2_out[6]
  PIN prt2_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.759 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4276 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 454.330000 0.000000 454.430000 0.520000 ;
    END
  END prt2_out[5]
  PIN prt2_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 540.130000 0.000000 540.230000 0.520000 ;
    END
  END prt2_out[4]
  PIN prt2_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.521 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3364 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 625.930000 0.000000 626.030000 0.520000 ;
    END
  END prt2_out[3]
  PIN prt2_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.783 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5332 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 711.730000 0.000000 711.830000 0.520000 ;
    END
  END prt2_out[2]
  PIN prt2_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.279 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2276 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 797.530000 0.000000 797.630000 0.520000 ;
    END
  END prt2_out[1]
  PIN prt2_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 883.330000 0.000000 883.430000 0.520000 ;
    END
  END prt2_out[0]
  PIN prt2_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.4635 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0394 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 293.325000 0.000000 293.425000 0.520000 ;
    END
  END prt2_dir[7]
  PIN prt2_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.7195 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2538 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 379.125000 0.000000 379.225000 0.520000 ;
    END
  END prt2_dir[6]
  PIN prt2_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1315 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.322 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2608 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 464.925000 0.000000 465.025000 0.520000 ;
    END
  END prt2_dir[5]
  PIN prt2_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3715 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6346 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 10.706 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.1504 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 550.725000 0.000000 550.825000 0.520000 ;
    END
  END prt2_dir[4]
  PIN prt2_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.5165 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3166 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 636.525000 0.000000 636.625000 0.520000 ;
    END
  END prt2_dir[3]
  PIN prt2_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4135 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8634 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 13.642 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.0688 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 722.325000 0.000000 722.425000 0.520000 ;
    END
  END prt2_dir[2]
  PIN prt2_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.3765 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6566 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 808.125000 0.000000 808.225000 0.520000 ;
    END
  END prt2_dir[1]
  PIN prt2_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.2785 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2254 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 893.925000 0.000000 894.025000 0.520000 ;
    END
  END prt2_dir[0]
  PIN prt2_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7035 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0954 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 8.922 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.3008 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 297.285000 0.000000 297.385000 0.520000 ;
    END
  END prt2_ren[7]
  PIN prt2_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.5435 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4794 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 383.085000 0.000000 383.185000 0.520000 ;
    END
  END prt2_ren[6]
  PIN prt2_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6945 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0558 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7808 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 468.885000 0.000000 468.985000 0.520000 ;
    END
  END prt2_ren[5]
  PIN prt2_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 11.562 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.9168 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 554.685000 0.000000 554.785000 0.520000 ;
    END
  END prt2_ren[4]
  PIN prt2_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4855 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1802 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.146 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2864 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 640.485000 0.000000 640.585000 0.520000 ;
    END
  END prt2_ren[3]
  PIN prt2_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6675 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.937 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.586 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4224 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 726.285000 0.000000 726.385000 0.520000 ;
    END
  END prt2_ren[2]
  PIN prt2_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.878 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5072 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 812.085000 0.000000 812.185000 0.520000 ;
    END
  END prt2_ren[1]
  PIN prt2_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.3095 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4058 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 897.885000 0.000000 897.985000 0.520000 ;
    END
  END prt2_ren[0]
  PIN prt3_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.5395 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 81.6618 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2  ;
    ANTENNAMAXAREACAR 537.19 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 2364.1 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 641.335000 0.520000 641.435000 ;
    END
  END prt3_in[7]
  PIN prt3_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4885 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.2374 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2  ;
    ANTENNAMAXAREACAR 573.146 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 2523.63 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 553.335000 0.520000 553.435000 ;
    END
  END prt3_in[6]
  PIN prt3_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4905 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0022 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 18.228 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.2912 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M3  ;
    ANTENNAMAXAREACAR 632.791 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 2787.4 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 1.89702 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 1.262 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5968 LAYER M4  ;
    ANTENNAGATEAREA 0.1038 LAYER M4  ;
    ANTENNAMAXAREACAR 644.949 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 2841.32 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.89702 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 465.335000 0.520000 465.435000 ;
    END
  END prt3_in[5]
  PIN prt3_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2925 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.287 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 3.602 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8928 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 14.706 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 64.7504 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M5  ;
    ANTENNAMAXAREACAR 150.916 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 666.035 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.19836 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 377.335000 0.520000 377.435000 ;
    END
  END prt3_in[4]
  PIN prt3_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1755 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7722 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 19.19 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.568 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 LAYER M3  ;
    ANTENNAMAXAREACAR 129.056 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 568.651 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 289.335000 0.520000 289.435000 ;
    END
  END prt3_in[3]
  PIN prt3_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0335 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9914 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 471.504 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 2078.03 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 201.335000 0.520000 201.435000 ;
    END
  END prt3_in[2]
  PIN prt3_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.5315 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.0266 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 4.258 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7792 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 459.769 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 2024.77 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 113.335000 0.520000 113.435000 ;
    END
  END prt3_in[1]
  PIN prt3_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8505 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1862 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 13.342 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.7488 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3  ;
    ANTENNAMAXAREACAR 409.205 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1783.97 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 25.335000 0.520000 25.435000 ;
    END
  END prt3_in[0]
  PIN prt3_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 14.903 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.6612 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 661.570000 0.520000 661.670000 ;
    END
  END prt3_out[7]
  PIN prt3_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 6.016 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.5584 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 573.570000 0.520000 573.670000 ;
    END
  END prt3_out[6]
  PIN prt3_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.036 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5584 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.726 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6384 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 485.570000 0.520000 485.670000 ;
    END
  END prt3_out[5]
  PIN prt3_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.137 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6468 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 397.570000 0.520000 397.670000 ;
    END
  END prt3_out[4]
  PIN prt3_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.615 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.394 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 309.570000 0.520000 309.670000 ;
    END
  END prt3_out[3]
  PIN prt3_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 9.4 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.448 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 221.570000 0.520000 221.670000 ;
    END
  END prt3_out[2]
  PIN prt3_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 13.25 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.344 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 133.570000 0.520000 133.670000 ;
    END
  END prt3_out[1]
  PIN prt3_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.959 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5076 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 45.570000 0.520000 45.670000 ;
    END
  END prt3_out[0]
  PIN prt3_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 13.8995 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.2458 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 650.975000 0.520000 651.075000 ;
    END
  END prt3_dir[7]
  PIN prt3_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.5686 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.786 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5024 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 562.975000 0.520000 563.075000 ;
    END
  END prt3_dir[6]
  PIN prt3_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 474.975000 0.520000 475.075000 ;
    END
  END prt3_dir[5]
  PIN prt3_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 15.562 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.5168 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 386.975000 0.520000 387.075000 ;
    END
  END prt3_dir[4]
  PIN prt3_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7515 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3066 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 16.766 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.8144 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.878 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9072 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 298.975000 0.520000 299.075000 ;
    END
  END prt3_dir[3]
  PIN prt3_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 14.7965 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.1486 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 210.975000 0.520000 211.075000 ;
    END
  END prt3_dir[2]
  PIN prt3_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 13.9165 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.3646 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 122.975000 0.520000 123.075000 ;
    END
  END prt3_dir[1]
  PIN prt3_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 2.8975 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.881 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 34.975000 0.520000 35.075000 ;
    END
  END prt3_dir[0]
  PIN prt3_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 14.2215 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.7066 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 647.015000 0.520000 647.115000 ;
    END
  END prt3_ren[7]
  PIN prt3_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6185 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.3654 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.166 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1744 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 559.015000 0.520000 559.115000 ;
    END
  END prt3_ren[6]
  PIN prt3_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.3862 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.042 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0288 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 471.015000 0.520000 471.115000 ;
    END
  END prt3_ren[5]
  PIN prt3_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4005 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7622 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 6.898 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.3952 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 383.015000 0.520000 383.115000 ;
    END
  END prt3_ren[4]
  PIN prt3_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2075 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.913 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 6.412 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3008 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 295.015000 0.520000 295.115000 ;
    END
  END prt3_ren[3]
  PIN prt3_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 7.1125 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.427 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 207.015000 0.520000 207.115000 ;
    END
  END prt3_ren[2]
  PIN prt3_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.1805 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.1942 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.506 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.8704 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 119.015000 0.520000 119.115000 ;
    END
  END prt3_ren[1]
  PIN prt3_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5805 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5542 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.4 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.048 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 0.000000 31.015000 0.520000 31.115000 ;
    END
  END prt3_ren[0]
  PIN prt4_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9642 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 25.812 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.661 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3  ;
    ANTENNAMAXAREACAR 412.374 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1807.8 LAYER M3  ;
    ANTENNAMAXCUTCAR 2.16802 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 646.165000 685.480000 646.265000 686.000000 ;
    END
  END prt4_in[7]
  PIN prt4_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9355 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5162 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 17.758 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.1792 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 5.078 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3872 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4  ;
    ANTENNAMAXAREACAR 67.1771 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 296.923 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 560.365000 685.480000 560.465000 686.000000 ;
    END
  END prt4_in[6]
  PIN prt4_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 7.602 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.4928 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 2.818 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4432 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4  ;
    ANTENNAMAXAREACAR 51.23 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 227.415 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.54769 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 474.565000 685.480000 474.665000 686.000000 ;
    END
  END prt4_in[5]
  PIN prt4_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7775 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.865 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M2  ;
    ANTENNAMAXAREACAR 184.919 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 814.374 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.186 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M3  ;
    ANTENNAGATEAREA 0.0369 LAYER M3  ;
    ANTENNAMAXAREACAR 189.959 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 837.745 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.622 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7808 LAYER M4  ;
    ANTENNAGATEAREA 0.1038 LAYER M4  ;
    ANTENNAMAXAREACAR 195.952 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 864.535 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 388.765000 685.480000 388.865000 686.000000 ;
    END
  END prt4_in[4]
  PIN prt4_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2485 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.9814 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M2  ;
    ANTENNAMAXAREACAR 203.121 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 892.851 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3  ;
    ANTENNAGATEAREA 0.1038 LAYER M3  ;
    ANTENNAMAXAREACAR 206.069 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 906.246 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 302.965000 685.480000 303.065000 686.000000 ;
    END
  END prt4_in[3]
  PIN prt4_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 12.94 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.024 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3  ;
    ANTENNAMAXAREACAR 290.29 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1277.85 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 217.165000 685.480000 217.265000 686.000000 ;
    END
  END prt4_in[2]
  PIN prt4_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.731 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 20.698 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.1152 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 6.598 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.0752 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4  ;
    ANTENNAMAXAREACAR 76.013 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 332.508 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.927362 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 131.365000 685.480000 131.465000 686.000000 ;
    END
  END prt4_in[1]
  PIN prt4_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2725 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 27.886 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.742 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3  ;
    ANTENNAMAXAREACAR 1077.86 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 4725.82 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 45.565000 685.480000 45.665000 686.000000 ;
    END
  END prt4_in[0]
  PIN prt4_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.652 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7766 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 47.6 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.536 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 625.930000 685.480000 626.030000 686.000000 ;
    END
  END prt4_out[7]
  PIN prt4_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.572 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4886 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 10.08 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.264 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 540.130000 685.480000 540.230000 686.000000 ;
    END
  END prt4_out[6]
  PIN prt4_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 13.922 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4902 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 454.330000 685.480000 454.430000 686.000000 ;
    END
  END prt4_out[5]
  PIN prt4_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.762 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5142 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 368.530000 685.480000 368.630000 686.000000 ;
    END
  END prt4_out[4]
  PIN prt4_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.968 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 6.038 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.6112 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 282.730000 685.480000 282.830000 686.000000 ;
    END
  END prt4_out[3]
  PIN prt4_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 14.342 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.1488 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 196.930000 685.480000 197.030000 686.000000 ;
    END
  END prt4_out[2]
  PIN prt4_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 111.130000 685.480000 111.230000 686.000000 ;
    END
  END prt4_out[1]
  PIN prt4_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 25.330000 685.480000 25.430000 686.000000 ;
    END
  END prt4_out[0]
  PIN prt4_dir[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 12.106 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.3104 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 636.525000 685.480000 636.625000 686.000000 ;
    END
  END prt4_dir[7]
  PIN prt4_dir[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.4965 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2286 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 550.725000 685.480000 550.825000 686.000000 ;
    END
  END prt4_dir[6]
  PIN prt4_dir[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.3005 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3222 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 464.925000 685.480000 465.025000 686.000000 ;
    END
  END prt4_dir[5]
  PIN prt4_dir[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.4995 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5978 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 379.125000 685.480000 379.225000 686.000000 ;
    END
  END prt4_dir[4]
  PIN prt4_dir[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.871 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8324 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.968 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.898 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5952 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 293.325000 685.480000 293.425000 686.000000 ;
    END
  END prt4_dir[3]
  PIN prt4_dir[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.491 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1604 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 13.522 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.5408 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 207.525000 685.480000 207.625000 686.000000 ;
    END
  END prt4_dir[2]
  PIN prt4_dir[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.722 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 73.6208 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 121.725000 685.480000 121.825000 686.000000 ;
    END
  END prt4_dir[1]
  PIN prt4_dir[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 35.925000 685.480000 36.025000 686.000000 ;
    END
  END prt4_dir[0]
  PIN prt4_ren[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5075 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.233 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 13.662 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.1568 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 640.485000 685.480000 640.585000 686.000000 ;
    END
  END prt4_ren[7]
  PIN prt4_ren[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.1385 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0534 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 554.685000 685.480000 554.785000 686.000000 ;
    END
  END prt4_ren[6]
  PIN prt4_ren[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2305 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4142 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 7.362 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.4368 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 468.885000 685.480000 468.985000 686.000000 ;
    END
  END prt4_ren[5]
  PIN prt4_ren[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.7205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5702 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 383.085000 685.480000 383.185000 686.000000 ;
    END
  END prt4_ren[4]
  PIN prt4_ren[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9985 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6374 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 297.285000 685.480000 297.385000 686.000000 ;
    END
  END prt4_ren[3]
  PIN prt4_ren[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6635 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9194 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 13.102 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.6928 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 211.485000 685.480000 211.585000 686.000000 ;
    END
  END prt4_ren[2]
  PIN prt4_ren[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8035 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5354 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 125.685000 685.480000 125.785000 686.000000 ;
    END
  END prt4_ren[1]
  PIN prt4_ren[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 16.762 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 73.7968 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 39.885000 685.480000 39.985000 686.000000 ;
    END
  END prt4_ren[0]
  PIN use_dac_glb_bias
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.7225 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.223 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 614.515000 399.000000 614.615000 ;
    END
  END use_dac_glb_bias
  PIN en_bias_buf
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.076 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.458 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0592 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 5.562 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 24.5168 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 11.078 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 48.7872 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 613.970000 399.000000 614.070000 ;
    END
  END en_bias_buf
  PIN en_bias_gen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.839 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1356 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.106 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.218 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4032 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 612.880000 399.000000 612.980000 ;
    END
  END en_bias_gen
  PIN BIAS_ADJ[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.843 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1972 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 609.610000 399.000000 609.710000 ;
    END
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 5.146 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6864 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 10.276 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 45.3024 LAYER M6  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6  ;
    ANTENNADIFFAREA 1.696 LAYER M7  ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M7  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M7  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M7  ;
    ANTENNAMAXAREACAR 171.894 LAYER M7  ;
    ANTENNAMAXSIDEAREACAR 758.69 LAYER M7  ;
    ANTENNAMAXCUTCAR 1.7316 LAYER VIA7  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 610.155000 399.000000 610.255000 ;
    END
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.998 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6352 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.818 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 43.2432 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6  ;
    ANTENNAMAXAREACAR 263.101 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1161.46 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 610.700000 399.000000 610.800000 ;
    END
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.002 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4528 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.158 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 2.186 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6624 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 11.058 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 48.6992 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6  ;
    ANTENNAMAXAREACAR 254.301 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1122.74 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.33333 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 611.245000 399.000000 611.345000 ;
    END
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5368 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.422 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3008 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 2.718 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0032 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.996 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 44.0704 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6  ;
    ANTENNAMAXAREACAR 242.482 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1070.52 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 611.790000 399.000000 611.890000 ;
    END
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.822 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0608 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 1.678 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4272 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.796 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 43.1904 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 612.335000 399.000000 612.435000 ;
    END
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.142 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.922 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7008 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 10.798 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 47.5552 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 601.980000 399.000000 602.080000 ;
    END
  END BIAS_DBP[13]
  PIN BIAS_DBP[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 5.166 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 22.7744 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 12.9 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 56.848 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6  ;
    ANTENNAMAXAREACAR 311.957 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1376.05 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 602.525000 399.000000 602.625000 ;
    END
  END BIAS_DBP[12]
  PIN BIAS_DBP[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.0816 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 5.566 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 24.5344 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 11.698 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 51.5152 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 603.070000 399.000000 603.170000 ;
    END
  END BIAS_DBP[11]
  PIN BIAS_DBP[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.692 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0255 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1562 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 603.615000 399.000000 603.715000 ;
    END
  END BIAS_DBP[10]
  PIN BIAS_DBP[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 5.002 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 22.0528 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 11.576 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 51.0224 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 604.160000 399.000000 604.260000 ;
    END
  END BIAS_DBP[9]
  PIN BIAS_DBP[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0675 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.341 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 604.705000 399.000000 604.805000 ;
    END
  END BIAS_DBP[8]
  PIN BIAS_DBP[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.847 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7268 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.662 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3568 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 605.250000 399.000000 605.350000 ;
    END
  END BIAS_DBP[7]
  PIN BIAS_DBP[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.164 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6096 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 605.795000 399.000000 605.895000 ;
    END
  END BIAS_DBP[6]
  PIN BIAS_DBP[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 4.456 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6944 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M6  ;
    ANTENNAMAXAREACAR 141.834 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 630.918 LAYER M6  ;
    ANTENNAMAXCUTCAR 2.18579 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 606.340000 399.000000 606.440000 ;
    END
  END BIAS_DBP[5]
  PIN BIAS_DBP[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.6585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9414 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 606.885000 399.000000 606.985000 ;
    END
  END BIAS_DBP[4]
  PIN BIAS_DBP[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.062 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3168 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 4.22 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.656 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 1.586 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0224 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 4.92 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6  ;
    ANTENNAMAXAREACAR 308.184 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1362.93 LAYER M6  ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 607.430000 399.000000 607.530000 ;
    END
  END BIAS_DBP[3]
  PIN BIAS_DBP[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.602 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0928 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 6.216 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 27.4384 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6  ;
    ANTENNAMAXAREACAR 240.482 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1065.04 LAYER M6  ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 607.975000 399.000000 608.075000 ;
    END
  END BIAS_DBP[2]
  PIN BIAS_DBP[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 608.520000 399.000000 608.620000 ;
    END
  END BIAS_DBP[1]
  PIN BIAS_DBP[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0885 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.856 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6544 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 2.726 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0384 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 5.578 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 24.5872 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6  ;
    ANTENNAMAXAREACAR 211.828 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 935.061 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 609.065000 399.000000 609.165000 ;
    END
  END BIAS_DBP[0]
  PIN BIAS_DBN[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 2.958 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0592 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 1.498 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6352 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 1.338 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9312 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 7.364 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 32.4896 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6  ;
    ANTENNAMAXAREACAR 119.773 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 529.356 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 579.090000 399.000000 579.190000 ;
    END
  END BIAS_DBN[13]
  PIN BIAS_DBN[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4055 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1842 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.086 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4224 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.968 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 4.738 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8912 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 579.635000 399.000000 579.735000 ;
    END
  END BIAS_DBN[12]
  PIN BIAS_DBN[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.597 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4268 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.968 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 4.002 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6528 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 580.180000 399.000000 580.280000 ;
    END
  END BIAS_DBN[11]
  PIN BIAS_DBN[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.968 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 5.538 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.4112 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 580.725000 399.000000 580.825000 ;
    END
  END BIAS_DBN[10]
  PIN BIAS_DBN[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.22 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.34 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 581.270000 399.000000 581.370000 ;
    END
  END BIAS_DBN[9]
  PIN BIAS_DBN[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.678 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0272 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 581.815000 399.000000 581.915000 ;
    END
  END BIAS_DBN[8]
  PIN BIAS_DBN[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.513 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3012 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.138 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 582.360000 399.000000 582.460000 ;
    END
  END BIAS_DBN[7]
  PIN BIAS_DBN[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4515 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0306 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.158 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 582.905000 399.000000 583.005000 ;
    END
  END BIAS_DBN[6]
  PIN BIAS_DBN[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 2.962 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0768 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.978 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 6.518 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 28.7232 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6  ;
    ANTENNAMAXAREACAR 356.214 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1572.49 LAYER M6  ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 583.450000 399.000000 583.550000 ;
    END
  END BIAS_DBN[5]
  PIN BIAS_DBN[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 2.498 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0352 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.506 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2704 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 7.278 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 32.0672 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER M6  ;
    ANTENNAMAXAREACAR 163.191 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 721.322 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.4245 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 583.995000 399.000000 584.095000 ;
    END
  END BIAS_DBN[4]
  PIN BIAS_DBN[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.833 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6652 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.766 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4144 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 584.540000 399.000000 584.640000 ;
    END
  END BIAS_DBN[3]
  PIN BIAS_DBN[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 5.282 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 23.2848 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.404 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 41.4656 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6  ;
    ANTENNAMAXAREACAR 210.85 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 929.492 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 585.085000 399.000000 585.185000 ;
    END
  END BIAS_DBN[2]
  PIN BIAS_DBN[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.822 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0608 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 4.362 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2368 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 7.874 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 34.7776 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6  ;
    ANTENNAMAXAREACAR 444.305 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1960.55 LAYER M6  ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 585.630000 399.000000 585.730000 ;
    END
  END BIAS_DBN[1]
  PIN BIAS_DBN[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 3.342 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7488 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.698 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1152 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 1.962 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6768 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.098 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 40.0752 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6  ;
    ANTENNAMAXAREACAR 260.281 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1148.84 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 586.175000 399.000000 586.275000 ;
    END
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 594.350000 399.000000 594.450000 ;
    END
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 594.895000 399.000000 594.995000 ;
    END
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.71 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.212 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 595.440000 399.000000 595.540000 ;
    END
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.3155 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4322 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 595.985000 399.000000 596.085000 ;
    END
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 596.530000 399.000000 596.630000 ;
    END
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2882 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 597.075000 399.000000 597.175000 ;
    END
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.0684 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 6.044 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.6816 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 4.642 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4688 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 7.622 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 33.5808 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6  ;
    ANTENNAMAXAREACAR 393.568 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1734.15 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 597.620000 399.000000 597.720000 ;
    END
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 1.506 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 13.234 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 58.3616 LAYER M6  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6  ;
    ANTENNADIFFAREA 1.696 LAYER M7  ;
    ANTENNAPARTIALMETALAREA 2.938 LAYER M7  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0592 LAYER M7  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7  ;
    ANTENNAMAXAREACAR 168.973 LAYER M7  ;
    ANTENNAMAXSIDEAREACAR 747.939 LAYER M7  ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA7  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 598.165000 399.000000 598.265000 ;
    END
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.958 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6592 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 598.710000 399.000000 598.810000 ;
    END
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.748 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3792 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 599.255000 399.000000 599.355000 ;
    END
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.142 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6248 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.548 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 599.800000 399.000000 599.900000 ;
    END
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 6.818 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0432 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4  ;
    ANTENNAMAXAREACAR 254.402 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 1119.75 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 600.345000 399.000000 600.445000 ;
    END
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.051 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2244 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.458 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.622 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7808 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 600.890000 399.000000 600.990000 ;
    END
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2445 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1198 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 2.562 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3168 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 4.138 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2512 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 2.832 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5928 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 4.564 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1696 LAYER M6  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6  ;
    ANTENNADIFFAREA 1.696 LAYER M7  ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M7  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M7  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7  ;
    ANTENNAMAXAREACAR 25.2836 LAYER M7  ;
    ANTENNAMAXSIDEAREACAR 114.411 LAYER M7  ;
    ANTENNAMAXCUTCAR 1.77994 LAYER VIA7  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 601.435000 399.000000 601.535000 ;
    END
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 3.318 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6432 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 4.922 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7008 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 1.062 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7168 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 4.522 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 19.9408 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6  ;
    ANTENNAMAXAREACAR 134.417 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 595.688 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 586.720000 399.000000 586.820000 ;
    END
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.502 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1264 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 2.478 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9472 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.086 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4224 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 5.338 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 23.5312 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6  ;
    ANTENNAMAXAREACAR 123.299 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 546.133 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 587.265000 399.000000 587.365000 ;
    END
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.358 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 2.878 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7072 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.968 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 3.538 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6112 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 587.810000 399.000000 587.910000 ;
    END
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 3.018 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3232 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 6.198 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 27.3152 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6  ;
    ANTENNAMAXAREACAR 96.1201 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 425.911 LAYER M6  ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 588.355000 399.000000 588.455000 ;
    END
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.422 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3008 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.118 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 40.1632 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6  ;
    ANTENNAMAXAREACAR 185.367 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 818.703 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 588.900000 399.000000 589.000000 ;
    END
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1415 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6666 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 2.862 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6368 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 6.618 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1632 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 2.618 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5632 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6  ;
    ANTENNAMAXAREACAR 105.601 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 467.73 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 589.445000 399.000000 589.545000 ;
    END
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4488 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 7.858 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.6192 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M5  ;
    ANTENNAMAXAREACAR 21.3408 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 90.5033 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 589.990000 399.000000 590.090000 ;
    END
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.418 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 7.176 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 31.6624 LAYER M6  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6  ;
    ANTENNADIFFAREA 1.696 LAYER M7  ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M7  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M7  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M7  ;
    ANTENNAMAXAREACAR 22.9342 LAYER M7  ;
    ANTENNAMAXSIDEAREACAR 104.73 LAYER M7  ;
    ANTENNAMAXCUTCAR 1.83333 LAYER VIA7  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 590.535000 399.000000 590.635000 ;
    END
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.326 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4784 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 9.142 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 40.3568 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6  ;
    ANTENNAMAXAREACAR 464.871 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 2053.54 LAYER M6  ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 591.080000 399.000000 591.180000 ;
    END
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.458 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 591.625000 399.000000 591.725000 ;
    END
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 6.978 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 30.7472 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M6  ;
    ANTENNAMAXAREACAR 187.406 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 815.547 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.64609 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 592.170000 399.000000 592.270000 ;
    END
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.982 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3648 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.158 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 2.386 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5424 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 7.318 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 32.2432 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 592.715000 399.000000 592.815000 ;
    END
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1012 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.482 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5648 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4112 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 1.742 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7088 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 6.916 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 30.5184 LAYER M6  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6  ;
    ANTENNADIFFAREA 1.696 LAYER M7  ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M7  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M7  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M7  ;
    ANTENNAMAXAREACAR 177.686 LAYER M7  ;
    ANTENNAMAXSIDEAREACAR 788.505 LAYER M7  ;
    ANTENNAMAXCUTCAR 3.55987 LAYER VIA7  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 593.260000 399.000000 593.360000 ;
    END
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0195 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.478 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1472 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 398.480000 593.805000 399.000000 593.905000 ;
    END
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.4835 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1714 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3  ;
    ANTENNAMAXAREACAR 11.8592 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 53.0667 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1047.865000 445.480000 1047.965000 446.000000 ;
    END
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.043 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5892 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.96 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 15.1 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 66.528 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M6  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6  ;
    ANTENNADIFFAREA 1.696 LAYER M7  ;
    ANTENNAPARTIALMETALAREA 5.392 LAYER M7  ;
    ANTENNAPARTIALMETALSIDEAREA 23.8128 LAYER M7  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0411 LAYER M7  ;
    ANTENNAMAXAREACAR 782.012 LAYER M7  ;
    ANTENNAMAXSIDEAREACAR 3436.03 LAYER M7  ;
    ANTENNAMAXCUTCAR 2.91971 LAYER VIA7  ;
    PORT
      LAYER M2 ;
        RECT 1048.410000 445.480000 1048.510000 446.000000 ;
    END
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6165 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7126 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1048.955000 445.480000 1049.055000 446.000000 ;
    END
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.493 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2132 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1049.500000 445.480000 1049.600000 446.000000 ;
    END
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3505 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5422 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.758 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3792 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3  ;
    ANTENNAMAXAREACAR 34.3916 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 152.317 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.323625 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1050.045000 445.480000 1050.145000 446.000000 ;
    END
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.241 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4604 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M2  ;
    ANTENNAMAXAREACAR 20.8803 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 91.4434 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.161812 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 1050.590000 445.480000 1050.690000 446.000000 ;
    END
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2505 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1022 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.488 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0352 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3  ;
    ANTENNAMAXAREACAR 44.7167 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 198.403 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1051.135000 445.480000 1051.235000 446.000000 ;
    END
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.224 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9856 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.802 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5728 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1051.680000 445.480000 1051.780000 446.000000 ;
    END
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3828 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.4995 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2418 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M4  ;
    ANTENNAMAXAREACAR 43.7167 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 194.737 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1052.225000 445.480000 1052.325000 446.000000 ;
    END
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.462 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4768 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3  ;
    ANTENNAMAXAREACAR 26.6833 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 118.323 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1052.770000 445.480000 1052.870000 446.000000 ;
    END
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1375 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.605 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.338 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9312 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4  ;
    ANTENNAMAXAREACAR 62.2091 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 274.036 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1053.315000 445.480000 1053.415000 446.000000 ;
    END
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.058 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7432 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.978 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3  ;
    ANTENNAMAXAREACAR 17.4009 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 77.3204 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.323625 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1053.860000 445.480000 1053.960000 446.000000 ;
    END
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1335 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5874 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 4.396 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4304 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1039.145000 445.480000 1039.245000 446.000000 ;
    END
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.511 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2484 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.486 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1824 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 7.118 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 31.3632 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1039.690000 445.480000 1039.790000 446.000000 ;
    END
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4695 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0658 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.5808 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1040.235000 445.480000 1040.335000 446.000000 ;
    END
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 5.258 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.1792 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1040.780000 445.480000 1040.880000 446.000000 ;
    END
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.071 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3124 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 2.438 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7712 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1041.325000 445.480000 1041.425000 446.000000 ;
    END
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.249 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0956 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.782 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6848 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1041.870000 445.480000 1041.970000 446.000000 ;
    END
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1042.415000 445.480000 1042.515000 446.000000 ;
    END
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.075 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.33 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 3.624 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0336 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M6  ;
    PORT
      LAYER M2 ;
        RECT 1042.960000 445.480000 1043.060000 446.000000 ;
    END
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.5295 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3298 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1043.505000 445.480000 1043.605000 446.000000 ;
    END
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.287 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6628 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.788 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3552 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.586 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 24.158 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 106.339 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M6  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6  ;
    ANTENNADIFFAREA 1.696 LAYER M7  ;
    ANTENNAPARTIALMETALAREA 2.602 LAYER M7  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4928 LAYER M7  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0481 LAYER M7  ;
    ANTENNAMAXAREACAR 279.371 LAYER M7  ;
    ANTENNAMAXSIDEAREACAR 1235.97 LAYER M7  ;
    ANTENNAMAXCUTCAR 2.2869 LAYER VIA7  ;
    PORT
      LAYER M2 ;
        RECT 1044.050000 445.480000 1044.150000 446.000000 ;
    END
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.4145 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8678 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1044.595000 445.480000 1044.695000 446.000000 ;
    END
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.466 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0944 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.058 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6992 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1045.140000 445.480000 1045.240000 446.000000 ;
    END
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.431 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8964 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.3785 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1094 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1045.685000 445.480000 1045.785000 446.000000 ;
    END
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.29 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.32 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1046.230000 445.480000 1046.330000 446.000000 ;
    END
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0915 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4026 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.342 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9488 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1046.775000 445.480000 1046.875000 446.000000 ;
    END
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6776 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.218 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4032 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1047.320000 445.480000 1047.420000 446.000000 ;
    END
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.602 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6928 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.598 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0752 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 607.010000 1139.520000 607.110000 ;
    END
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.378 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1072 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 607.555000 1139.520000 607.655000 ;
    END
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.742 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3088 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 608.100000 1139.520000 608.200000 ;
    END
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.058 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6992 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 608.645000 1139.520000 608.745000 ;
    END
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 2.358 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3752 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 609.190000 1139.520000 609.290000 ;
    END
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.3705 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0742 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 609.735000 1139.520000 609.835000 ;
    END
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.106 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 610.280000 1139.520000 610.380000 ;
    END
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.906 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0304 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 610.825000 1139.520000 610.925000 ;
    END
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.217 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9988 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 611.370000 1139.520000 611.470000 ;
    END
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0305 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1342 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.502 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 611.915000 1139.520000 612.015000 ;
    END
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.068 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.726 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2384 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 612.460000 1139.520000 612.560000 ;
    END
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0195 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.818 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6432 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 613.005000 1139.520000 613.105000 ;
    END
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.074 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3256 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 613.550000 1139.520000 613.650000 ;
    END
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0845 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4158 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 614.095000 1139.520000 614.195000 ;
    END
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5375 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.409 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2  ;
    ANTENNAMAXAREACAR 9.87374 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 42.2164 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3  ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 13.6544 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 59.4863 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.978 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M4  ;
    ANTENNAGATEAREA 0.0693 LAYER M4  ;
    ANTENNAMAXAREACAR 27.767 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 122.216 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1029.335000 445.480000 1029.435000 446.000000 ;
    END
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 2.498 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9912 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 29.816 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 131.278 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5  ;
    ANTENNADIFFAREA 1.696 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 6.166 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 27.1744 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6  ;
    ANTENNAMAXAREACAR 390.539 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 1721.21 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 1029.880000 445.480000 1029.980000 446.000000 ;
    END
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.5105 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2902 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1030.425000 445.480000 1030.525000 446.000000 ;
    END
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.379 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0676 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2  ;
    ANTENNAMAXAREACAR 20.8189 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 90.3867 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.446 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0064 LAYER M3  ;
    ANTENNAGATEAREA 0.0693 LAYER M3  ;
    ANTENNAMAXAREACAR 27.2547 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 119.339 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1030.970000 445.480000 1031.070000 446.000000 ;
    END
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7975 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.509 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.886 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9424 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1031.515000 445.480000 1031.615000 446.000000 ;
    END
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.888 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9512 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1032.060000 445.480000 1032.160000 446.000000 ;
    END
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1115 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4906 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.658 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9392 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4  ;
    ANTENNAMAXAREACAR 122.506 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 538.984 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1032.605000 445.480000 1032.705000 446.000000 ;
    END
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.551 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4244 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.432 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.582 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6048 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 1.558 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5  ;
    ANTENNAMAXAREACAR 49.4664 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 214.252 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1033.150000 445.480000 1033.250000 446.000000 ;
    END
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1225 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.1424 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7696 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 3.218 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2032 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5  ;
    ANTENNAMAXAREACAR 64.3912 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 285.502 LAYER M5  ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1033.695000 445.480000 1033.795000 446.000000 ;
    END
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.047 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.142 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0688 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 2.942 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9888 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5  ;
    ANTENNAMAXAREACAR 79.0376 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 347.744 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1034.240000 445.480000 1034.340000 446.000000 ;
    END
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1775 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.781 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1034.785000 445.480000 1034.885000 446.000000 ;
    END
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.391 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7204 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.502 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1035.330000 445.480000 1035.430000 446.000000 ;
    END
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.4885 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1494 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1026.065000 445.480000 1026.165000 446.000000 ;
    END
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.107 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8708 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.896 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8304 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3  ;
    ANTENNAMAXAREACAR 48.9806 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 217.107 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1026.610000 445.480000 1026.710000 446.000000 ;
    END
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.371 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6324 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.138 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.1 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.928 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 2.286 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1024 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5  ;
    ANTENNAMAXAREACAR 55.6214 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 247.152 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 1027.155000 445.480000 1027.255000 446.000000 ;
    END
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.129 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5676 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.958 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4  ;
    ANTENNAMAXAREACAR 79.1489 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 349.961 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.809061 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 1027.700000 445.480000 1027.800000 446.000000 ;
    END
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1665 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7326 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1028.245000 445.480000 1028.345000 446.000000 ;
    END
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.685 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.014 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.438 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9712 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1028.790000 445.480000 1028.890000 446.000000 ;
    END
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7015 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0866 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.858 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8192 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1022.795000 445.480000 1022.895000 446.000000 ;
    END
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.696 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.19 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.48 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 LAYER M3  ;
    ANTENNAMAXAREACAR 95.7067 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 421.249 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.666667 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1023.340000 445.480000 1023.440000 446.000000 ;
    END
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.553 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4772 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1023.885000 445.480000 1023.985000 446.000000 ;
    END
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.385 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.694 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.898 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9952 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1024.430000 445.480000 1024.530000 446.000000 ;
    END
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6195 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7258 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.418 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2832 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1024.975000 445.480000 1025.075000 446.000000 ;
    END
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.24 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1025.520000 445.480000 1025.620000 446.000000 ;
    END
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.993 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.0572 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 599.380000 1139.520000 599.480000 ;
    END
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.698 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1152 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 599.925000 1139.520000 600.025000 ;
    END
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.22 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.948 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 600.470000 1139.520000 600.570000 ;
    END
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.278 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6672 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 601.015000 1139.520000 601.115000 ;
    END
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.818 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6432 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 601.560000 1139.520000 601.660000 ;
    END
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.142 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 602.105000 1139.520000 602.205000 ;
    END
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.082 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8048 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 602.650000 1139.520000 602.750000 ;
    END
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 603.195000 1139.520000 603.295000 ;
    END
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.344 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6016 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 603.740000 1139.520000 603.840000 ;
    END
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.3295 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4938 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 1.298 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7552 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 604.285000 1139.520000 604.385000 ;
    END
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 604.830000 1139.520000 604.930000 ;
    END
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.622 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7808 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 605.375000 1139.520000 605.475000 ;
    END
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.308 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 605.920000 1139.520000 606.020000 ;
    END
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.0275 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.165 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1139.000000 606.465000 1139.520000 606.565000 ;
    END
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.186 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8184 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 13.142 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.8688 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3  ;
    ANTENNAMAXAREACAR 341.62 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1504.42 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.755668 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 1008.030000 445.480000 1008.130000 446.000000 ;
    END
  END dsadc_conv_done
  PIN dsadc_en
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.237 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0868 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.682 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0448 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 5.804 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 25.6256 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1038.600000 445.480000 1038.700000 446.000000 ;
    END
  END dsadc_en
  PIN dsadc_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 9.224 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3224 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1037.510000 445.480000 1037.610000 446.000000 ;
    END
  END dsadc_clk
  PIN dsadc_switch[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.111 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4884 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.1205 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5742 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1035.875000 445.480000 1035.975000 446.000000 ;
    END
  END dsadc_switch[2]
  PIN dsadc_switch[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.584 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5696 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.618 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1632 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1036.420000 445.480000 1036.520000 446.000000 ;
    END
  END dsadc_switch[1]
  PIN dsadc_switch[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.291 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2804 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1036.965000 445.480000 1037.065000 446.000000 ;
    END
  END dsadc_switch[0]
  PIN dac_en_pot
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1665 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7326 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNADIFFAREA 1.696 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 5.198 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9152 LAYER M5  ;
    PORT
      LAYER M2 ;
        RECT 1038.055000 445.480000 1038.155000 446.000000 ;
    END
  END dac_en_pot
  PIN adc_ext_in
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.571 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5124 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 4.198 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.5152 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1022.250000 445.480000 1022.350000 446.000000 ;
    END
  END adc_ext_in
  PIN atp_en
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.462 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4768 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNADIFFAREA 1.696 LAYER M4  ;
    ANTENNAPARTIALMETALAREA 0.562 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5168 LAYER M4  ;
    PORT
      LAYER M2 ;
        RECT 1020.615000 445.480000 1020.715000 446.000000 ;
    END
  END atp_en
  PIN atp_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.364 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6456 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 1021.160000 445.480000 1021.260000 446.000000 ;
    END
  END atp_sel
  PIN adc_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3095 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3618 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 3.922 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.3008 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 1021.705000 445.480000 1021.805000 446.000000 ;
    END
  END adc_sel
  PIN saradc_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNADIFFAREA 1.696 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 65.902 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.6682 LAYER M3  ;
    PORT
      LAYER M2 ;
        RECT 884.605000 445.480000 884.705000 446.000000 ;
    END
  END saradc_clk
  PIN saradc_rdy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.481 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2484 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2  ;
    ANTENNAMAXAREACAR 25.5908 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 110.807 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2  ;
    PORT
      LAYER M2 ;
        RECT 884.205000 445.480000 884.305000 446.000000 ;
    END
  END saradc_rdy
  PIN saradc_rst
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.696 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.291 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2804 LAYER M2  ;
    PORT
      LAYER M2 ;
        RECT 883.805000 445.480000 883.905000 446.000000 ;
    END
  END saradc_rst
  PIN saradc_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8825 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.883 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 9.402 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.4128 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3  ;
    ANTENNAMAXAREACAR 272.166 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1190.89 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 883.405000 445.480000 883.505000 446.000000 ;
    END
  END saradc_data[9]
  PIN saradc_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4055 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8282 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 6.378 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.1072 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M4  ;
    ANTENNAMAXAREACAR 47.5642 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 211.683 LAYER M4  ;
    ANTENNAMAXCUTCAR 1.25945 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 883.005000 445.480000 883.105000 446.000000 ;
    END
  END saradc_data[8]
  PIN saradc_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4315 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8986 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 10.482 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.1648 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3  ;
    ANTENNAMAXAREACAR 279.37 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1226.55 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 882.605000 445.480000 882.705000 446.000000 ;
    END
  END saradc_data[7]
  PIN saradc_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.271 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1924 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 11.1335 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.0314 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3  ;
    ANTENNAMAXAREACAR 290.249 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1267.37 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 882.205000 445.480000 882.305000 446.000000 ;
    END
  END saradc_data[6]
  PIN saradc_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6755 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9722 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.098 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8752 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.266 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 12.638 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 55.6512 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 1.358 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0192 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M6  ;
    ANTENNAMAXAREACAR 125.013 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 547.259 LAYER M6  ;
    ANTENNAMAXCUTCAR 2.51889 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 881.805000 445.480000 881.905000 446.000000 ;
    END
  END saradc_data[5]
  PIN saradc_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5465 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4046 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 9.158 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.3392 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3  ;
    ANTENNAMAXAREACAR 246.725 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1083.64 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 881.405000 445.480000 881.505000 446.000000 ;
    END
  END saradc_data[4]
  PIN saradc_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1825 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.803 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.522 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7408 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 9.818 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 43.2432 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5  ;
    ANTENNAMAXAREACAR 342.393 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1508.99 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.01511 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 881.005000 445.480000 881.105000 446.000000 ;
    END
  END saradc_data[3]
  PIN saradc_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6425 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.827 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 11.258 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.5792 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3  ;
    ANTENNAMAXAREACAR 304.861 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 1338.35 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 880.605000 445.480000 880.705000 446.000000 ;
    END
  END saradc_data[2]
  PIN saradc_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.171 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7524 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.3135 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8234 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.606 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7104 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 9.938 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 43.7712 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5  ;
    ANTENNAMAXAREACAR 390.453 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1721.18 LAYER M5  ;
    ANTENNAMAXCUTCAR 2.01511 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 880.205000 445.480000 880.305000 446.000000 ;
    END
  END saradc_data[1]
  PIN saradc_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0395 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1738 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.566 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5344 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 13.678 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 60.2272 LAYER M5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5  ;
    ANTENNAMAXAREACAR 419.27 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 1846.5 LAYER M5  ;
    ANTENNAMAXCUTCAR 1.76322 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 879.805000 445.480000 879.905000 446.000000 ;
    END
  END saradc_data[0]
  PIN a0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[31]
  PIN a0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[30]
  PIN a0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[29]
  PIN a0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[28]
  PIN a0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[27]
  PIN a0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[26]
  PIN a0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[25]
  PIN a0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[24]
  PIN a0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[23]
  PIN a0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[22]
  PIN a0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[21]
  PIN a0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[20]
  PIN a0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[19]
  PIN a0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[18]
  PIN a0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[17]
  PIN a0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[16]
  PIN a0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[15]
  PIN a0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[14]
  PIN a0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[13]
  PIN a0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[12]
  PIN a0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[11]
  PIN a0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[10]
  PIN a0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[9]
  PIN a0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[8]
  PIN a0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[7]
  PIN a0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[6]
  PIN a0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[5]
  PIN a0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[4]
  PIN a0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[3]
  PIN a0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[2]
  PIN a0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[1]
  PIN a0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END a0[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M7 ;
        RECT 51.000000 0.000000 56.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 51.000000 681.000000 56.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 101.000000 0.000000 106.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 101.000000 681.000000 106.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 151.000000 0.000000 156.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 151.000000 681.000000 156.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 201.000000 0.000000 206.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 201.000000 681.000000 206.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 251.000000 0.000000 256.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 251.000000 681.000000 256.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 301.000000 0.000000 306.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 301.000000 681.000000 306.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 351.000000 0.000000 356.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 351.000000 681.000000 356.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 0.000000 406.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 501.000000 406.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 656.000000 406.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 401.000000 681.000000 406.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 0.000000 456.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 501.000000 456.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 656.000000 456.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 451.000000 681.000000 456.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 0.000000 506.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 501.000000 506.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 656.000000 506.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 501.000000 681.000000 506.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 0.000000 556.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 501.000000 556.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 656.000000 556.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 551.000000 681.000000 556.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 0.000000 606.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 501.000000 606.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 656.000000 606.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 601.000000 681.000000 606.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 0.000000 656.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 501.000000 656.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 656.000000 656.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 651.000000 681.000000 656.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 701.000000 0.000000 706.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 701.000000 501.000000 706.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 751.000000 0.000000 756.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 751.000000 441.000000 756.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 801.000000 0.000000 806.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 801.000000 441.000000 806.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 851.000000 0.000000 856.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 851.000000 441.000000 856.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 901.000000 0.000000 906.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 901.000000 441.000000 906.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 951.000000 0.000000 956.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 951.000000 441.000000 956.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1001.000000 0.000000 1006.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1001.000000 441.000000 1006.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1051.000000 0.000000 1056.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1051.000000 441.000000 1056.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1101.000000 0.000000 1106.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1101.000000 441.000000 1106.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1151.000000 0.000000 1156.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1151.000000 681.000000 1156.000000 686.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER M2 ;
        RECT 4.000000 5.850000 14.000000 6.150000 ;
        RECT 51.000000 5.850000 56.000000 6.150000 ;
        RECT 51.000000 1.850000 56.000000 2.150000 ;
        RECT 101.000000 1.850000 106.000000 2.150000 ;
        RECT 101.000000 5.850000 106.000000 6.150000 ;
        RECT 151.000000 1.850000 156.000000 2.150000 ;
        RECT 151.000000 5.850000 156.000000 6.150000 ;
        RECT 201.000000 1.850000 206.000000 2.150000 ;
        RECT 201.000000 5.850000 206.000000 6.150000 ;
        RECT 251.000000 1.850000 256.000000 2.150000 ;
        RECT 251.000000 5.850000 256.000000 6.150000 ;
        RECT 301.000000 1.850000 306.000000 2.150000 ;
        RECT 301.000000 5.850000 306.000000 6.150000 ;
        RECT 351.000000 1.850000 356.000000 2.150000 ;
        RECT 351.000000 5.850000 356.000000 6.150000 ;
        RECT 401.000000 1.850000 406.000000 2.150000 ;
        RECT 401.000000 5.850000 406.000000 6.150000 ;
        RECT 451.000000 1.850000 456.000000 2.150000 ;
        RECT 451.000000 5.850000 456.000000 6.150000 ;
        RECT 501.000000 1.850000 506.000000 2.150000 ;
        RECT 501.000000 5.850000 506.000000 6.150000 ;
        RECT 551.000000 1.850000 556.000000 2.150000 ;
        RECT 551.000000 5.850000 556.000000 6.150000 ;
        RECT 4.000000 265.850000 14.000000 266.150000 ;
        RECT 4.000000 261.850000 14.000000 262.150000 ;
        RECT 51.000000 265.850000 56.000000 266.150000 ;
        RECT 51.000000 261.850000 56.000000 262.150000 ;
        RECT 101.000000 265.850000 106.000000 266.150000 ;
        RECT 101.000000 261.850000 106.000000 262.150000 ;
        RECT 51.000000 305.850000 56.000000 306.150000 ;
        RECT 4.000000 305.850000 14.000000 306.150000 ;
        RECT 4.000000 285.850000 14.000000 286.150000 ;
        RECT 4.000000 281.850000 14.000000 282.150000 ;
        RECT 4.000000 269.850000 14.000000 270.150000 ;
        RECT 4.000000 273.850000 14.000000 274.150000 ;
        RECT 4.000000 277.850000 14.000000 278.150000 ;
        RECT 4.000000 289.850000 14.000000 290.150000 ;
        RECT 4.000000 293.850000 14.000000 294.150000 ;
        RECT 4.000000 297.850000 14.000000 298.150000 ;
        RECT 4.000000 301.850000 14.000000 302.150000 ;
        RECT 51.000000 269.850000 56.000000 270.150000 ;
        RECT 51.000000 273.850000 56.000000 274.150000 ;
        RECT 51.000000 277.850000 56.000000 278.150000 ;
        RECT 51.000000 281.850000 56.000000 282.150000 ;
        RECT 51.000000 285.850000 56.000000 286.150000 ;
        RECT 51.000000 301.850000 56.000000 302.150000 ;
        RECT 51.000000 297.850000 56.000000 298.150000 ;
        RECT 51.000000 293.850000 56.000000 294.150000 ;
        RECT 51.000000 289.850000 56.000000 290.150000 ;
        RECT 4.000000 321.850000 14.000000 322.150000 ;
        RECT 4.000000 317.850000 14.000000 318.150000 ;
        RECT 4.000000 309.850000 14.000000 310.150000 ;
        RECT 4.000000 313.850000 14.000000 314.150000 ;
        RECT 4.000000 325.850000 14.000000 326.150000 ;
        RECT 4.000000 329.850000 14.000000 330.150000 ;
        RECT 4.000000 333.850000 14.000000 334.150000 ;
        RECT 4.000000 337.850000 14.000000 338.150000 ;
        RECT 4.000000 341.850000 14.000000 342.150000 ;
        RECT 51.000000 313.850000 56.000000 314.150000 ;
        RECT 51.000000 309.850000 56.000000 310.150000 ;
        RECT 51.000000 317.850000 56.000000 318.150000 ;
        RECT 51.000000 321.850000 56.000000 322.150000 ;
        RECT 51.000000 341.850000 56.000000 342.150000 ;
        RECT 51.000000 337.850000 56.000000 338.150000 ;
        RECT 51.000000 333.850000 56.000000 334.150000 ;
        RECT 51.000000 329.850000 56.000000 330.150000 ;
        RECT 51.000000 325.850000 56.000000 326.150000 ;
        RECT 101.000000 305.850000 106.000000 306.150000 ;
        RECT 101.000000 285.850000 106.000000 286.150000 ;
        RECT 101.000000 269.850000 106.000000 270.150000 ;
        RECT 101.000000 273.850000 106.000000 274.150000 ;
        RECT 101.000000 277.850000 106.000000 278.150000 ;
        RECT 101.000000 281.850000 106.000000 282.150000 ;
        RECT 101.000000 301.850000 106.000000 302.150000 ;
        RECT 101.000000 297.850000 106.000000 298.150000 ;
        RECT 101.000000 293.850000 106.000000 294.150000 ;
        RECT 101.000000 289.850000 106.000000 290.150000 ;
        RECT 101.000000 321.850000 106.000000 322.150000 ;
        RECT 101.000000 317.850000 106.000000 318.150000 ;
        RECT 101.000000 313.850000 106.000000 314.150000 ;
        RECT 101.000000 309.850000 106.000000 310.150000 ;
        RECT 101.000000 325.850000 106.000000 326.150000 ;
        RECT 101.000000 329.850000 106.000000 330.150000 ;
        RECT 101.000000 333.850000 106.000000 334.150000 ;
        RECT 101.000000 337.850000 106.000000 338.150000 ;
        RECT 101.000000 341.850000 106.000000 342.150000 ;
        RECT 151.000000 261.850000 156.000000 262.150000 ;
        RECT 151.000000 265.850000 156.000000 266.150000 ;
        RECT 201.000000 265.850000 206.000000 266.150000 ;
        RECT 201.000000 261.850000 206.000000 262.150000 ;
        RECT 251.000000 265.850000 256.000000 266.150000 ;
        RECT 251.000000 261.850000 256.000000 262.150000 ;
        RECT 201.000000 305.850000 206.000000 306.150000 ;
        RECT 151.000000 305.850000 156.000000 306.150000 ;
        RECT 151.000000 277.850000 156.000000 278.150000 ;
        RECT 151.000000 273.850000 156.000000 274.150000 ;
        RECT 151.000000 269.850000 156.000000 270.150000 ;
        RECT 151.000000 281.850000 156.000000 282.150000 ;
        RECT 151.000000 285.850000 156.000000 286.150000 ;
        RECT 151.000000 289.850000 156.000000 290.150000 ;
        RECT 151.000000 293.850000 156.000000 294.150000 ;
        RECT 151.000000 297.850000 156.000000 298.150000 ;
        RECT 151.000000 301.850000 156.000000 302.150000 ;
        RECT 201.000000 269.850000 206.000000 270.150000 ;
        RECT 201.000000 273.850000 206.000000 274.150000 ;
        RECT 201.000000 277.850000 206.000000 278.150000 ;
        RECT 201.000000 281.850000 206.000000 282.150000 ;
        RECT 201.000000 285.850000 206.000000 286.150000 ;
        RECT 201.000000 301.850000 206.000000 302.150000 ;
        RECT 201.000000 297.850000 206.000000 298.150000 ;
        RECT 201.000000 293.850000 206.000000 294.150000 ;
        RECT 201.000000 289.850000 206.000000 290.150000 ;
        RECT 151.000000 313.850000 156.000000 314.150000 ;
        RECT 151.000000 309.850000 156.000000 310.150000 ;
        RECT 151.000000 321.850000 156.000000 322.150000 ;
        RECT 151.000000 317.850000 156.000000 318.150000 ;
        RECT 151.000000 329.850000 156.000000 330.150000 ;
        RECT 151.000000 325.850000 156.000000 326.150000 ;
        RECT 151.000000 333.850000 156.000000 334.150000 ;
        RECT 151.000000 337.850000 156.000000 338.150000 ;
        RECT 151.000000 341.850000 156.000000 342.150000 ;
        RECT 201.000000 313.850000 206.000000 314.150000 ;
        RECT 201.000000 309.850000 206.000000 310.150000 ;
        RECT 201.000000 317.850000 206.000000 318.150000 ;
        RECT 201.000000 321.850000 206.000000 322.150000 ;
        RECT 201.000000 341.850000 206.000000 342.150000 ;
        RECT 201.000000 337.850000 206.000000 338.150000 ;
        RECT 201.000000 333.850000 206.000000 334.150000 ;
        RECT 201.000000 329.850000 206.000000 330.150000 ;
        RECT 201.000000 325.850000 206.000000 326.150000 ;
        RECT 251.000000 305.850000 256.000000 306.150000 ;
        RECT 251.000000 285.850000 256.000000 286.150000 ;
        RECT 251.000000 269.850000 256.000000 270.150000 ;
        RECT 251.000000 273.850000 256.000000 274.150000 ;
        RECT 251.000000 277.850000 256.000000 278.150000 ;
        RECT 251.000000 281.850000 256.000000 282.150000 ;
        RECT 251.000000 293.850000 256.000000 294.150000 ;
        RECT 251.000000 289.850000 256.000000 290.150000 ;
        RECT 251.000000 301.850000 256.000000 302.150000 ;
        RECT 251.000000 297.850000 256.000000 298.150000 ;
        RECT 251.000000 321.850000 256.000000 322.150000 ;
        RECT 251.000000 317.850000 256.000000 318.150000 ;
        RECT 251.000000 313.850000 256.000000 314.150000 ;
        RECT 251.000000 309.850000 256.000000 310.150000 ;
        RECT 251.000000 325.850000 256.000000 326.150000 ;
        RECT 251.000000 329.850000 256.000000 330.150000 ;
        RECT 251.000000 337.850000 256.000000 338.150000 ;
        RECT 251.000000 333.850000 256.000000 334.150000 ;
        RECT 251.000000 341.850000 256.000000 342.150000 ;
        RECT 301.000000 265.850000 306.000000 266.150000 ;
        RECT 301.000000 261.850000 306.000000 262.150000 ;
        RECT 351.000000 265.850000 356.000000 266.150000 ;
        RECT 351.000000 261.850000 356.000000 262.150000 ;
        RECT 401.000000 261.850000 406.000000 262.150000 ;
        RECT 401.000000 265.850000 406.000000 266.150000 ;
        RECT 351.000000 305.850000 356.000000 306.150000 ;
        RECT 301.000000 305.850000 306.000000 306.150000 ;
        RECT 301.000000 277.850000 306.000000 278.150000 ;
        RECT 301.000000 269.850000 306.000000 270.150000 ;
        RECT 301.000000 273.850000 306.000000 274.150000 ;
        RECT 301.000000 281.850000 306.000000 282.150000 ;
        RECT 301.000000 285.850000 306.000000 286.150000 ;
        RECT 301.000000 293.850000 306.000000 294.150000 ;
        RECT 301.000000 289.850000 306.000000 290.150000 ;
        RECT 301.000000 301.850000 306.000000 302.150000 ;
        RECT 301.000000 297.850000 306.000000 298.150000 ;
        RECT 351.000000 269.850000 356.000000 270.150000 ;
        RECT 351.000000 273.850000 356.000000 274.150000 ;
        RECT 351.000000 277.850000 356.000000 278.150000 ;
        RECT 351.000000 281.850000 356.000000 282.150000 ;
        RECT 351.000000 285.850000 356.000000 286.150000 ;
        RECT 351.000000 301.850000 356.000000 302.150000 ;
        RECT 351.000000 297.850000 356.000000 298.150000 ;
        RECT 351.000000 293.850000 356.000000 294.150000 ;
        RECT 351.000000 289.850000 356.000000 290.150000 ;
        RECT 301.000000 313.850000 306.000000 314.150000 ;
        RECT 301.000000 309.850000 306.000000 310.150000 ;
        RECT 301.000000 317.850000 306.000000 318.150000 ;
        RECT 301.000000 321.850000 306.000000 322.150000 ;
        RECT 301.000000 329.850000 306.000000 330.150000 ;
        RECT 301.000000 325.850000 306.000000 326.150000 ;
        RECT 301.000000 341.850000 306.000000 342.150000 ;
        RECT 301.000000 337.850000 306.000000 338.150000 ;
        RECT 301.000000 333.850000 306.000000 334.150000 ;
        RECT 351.000000 313.850000 356.000000 314.150000 ;
        RECT 351.000000 309.850000 356.000000 310.150000 ;
        RECT 351.000000 317.850000 356.000000 318.150000 ;
        RECT 351.000000 321.850000 356.000000 322.150000 ;
        RECT 351.000000 341.850000 356.000000 342.150000 ;
        RECT 351.000000 337.850000 356.000000 338.150000 ;
        RECT 351.000000 333.850000 356.000000 334.150000 ;
        RECT 351.000000 329.850000 356.000000 330.150000 ;
        RECT 351.000000 325.850000 356.000000 326.150000 ;
        RECT 401.000000 305.850000 406.000000 306.150000 ;
        RECT 401.000000 277.850000 406.000000 278.150000 ;
        RECT 401.000000 269.850000 406.000000 270.150000 ;
        RECT 401.000000 273.850000 406.000000 274.150000 ;
        RECT 401.000000 285.850000 406.000000 286.150000 ;
        RECT 401.000000 281.850000 406.000000 282.150000 ;
        RECT 401.000000 301.850000 406.000000 302.150000 ;
        RECT 401.000000 297.850000 406.000000 298.150000 ;
        RECT 401.000000 293.850000 406.000000 294.150000 ;
        RECT 401.000000 289.850000 406.000000 290.150000 ;
        RECT 401.000000 313.850000 406.000000 314.150000 ;
        RECT 401.000000 309.850000 406.000000 310.150000 ;
        RECT 401.000000 317.850000 406.000000 318.150000 ;
        RECT 401.000000 321.850000 406.000000 322.150000 ;
        RECT 401.000000 329.850000 406.000000 330.150000 ;
        RECT 401.000000 325.850000 406.000000 326.150000 ;
        RECT 401.000000 333.850000 406.000000 334.150000 ;
        RECT 401.000000 337.850000 406.000000 338.150000 ;
        RECT 401.000000 341.850000 406.000000 342.150000 ;
        RECT 451.000000 265.850000 456.000000 266.150000 ;
        RECT 451.000000 261.850000 456.000000 262.150000 ;
        RECT 501.000000 261.850000 506.000000 262.150000 ;
        RECT 501.000000 265.850000 506.000000 266.150000 ;
        RECT 551.000000 265.850000 556.000000 266.150000 ;
        RECT 551.000000 261.850000 556.000000 262.150000 ;
        RECT 501.000000 305.850000 506.000000 306.150000 ;
        RECT 451.000000 277.850000 456.000000 278.150000 ;
        RECT 451.000000 273.850000 456.000000 274.150000 ;
        RECT 451.000000 269.850000 456.000000 270.150000 ;
        RECT 451.000000 285.850000 456.000000 286.150000 ;
        RECT 451.000000 281.850000 456.000000 282.150000 ;
        RECT 451.000000 293.850000 456.000000 294.150000 ;
        RECT 451.000000 289.850000 456.000000 290.150000 ;
        RECT 451.000000 297.850000 456.000000 298.150000 ;
        RECT 501.000000 277.850000 506.000000 278.150000 ;
        RECT 501.000000 269.850000 506.000000 270.150000 ;
        RECT 501.000000 273.850000 506.000000 274.150000 ;
        RECT 501.000000 281.850000 506.000000 282.150000 ;
        RECT 501.000000 285.850000 506.000000 286.150000 ;
        RECT 501.000000 289.850000 506.000000 290.150000 ;
        RECT 501.000000 293.850000 506.000000 294.150000 ;
        RECT 501.000000 297.850000 506.000000 298.150000 ;
        RECT 501.000000 301.850000 506.000000 302.150000 ;
        RECT 451.000000 321.850000 456.000000 322.150000 ;
        RECT 451.000000 333.850000 456.000000 334.150000 ;
        RECT 451.000000 329.850000 456.000000 330.150000 ;
        RECT 451.000000 325.850000 456.000000 326.150000 ;
        RECT 451.000000 337.850000 456.000000 338.150000 ;
        RECT 451.000000 341.850000 456.000000 342.150000 ;
        RECT 501.000000 313.850000 506.000000 314.150000 ;
        RECT 501.000000 309.850000 506.000000 310.150000 ;
        RECT 501.000000 317.850000 506.000000 318.150000 ;
        RECT 501.000000 321.850000 506.000000 322.150000 ;
        RECT 501.000000 329.850000 506.000000 330.150000 ;
        RECT 501.000000 325.850000 506.000000 326.150000 ;
        RECT 501.000000 333.850000 506.000000 334.150000 ;
        RECT 501.000000 337.850000 506.000000 338.150000 ;
        RECT 501.000000 341.850000 506.000000 342.150000 ;
        RECT 551.000000 305.850000 556.000000 306.150000 ;
        RECT 551.000000 281.850000 556.000000 282.150000 ;
        RECT 551.000000 277.850000 556.000000 278.150000 ;
        RECT 551.000000 273.850000 556.000000 274.150000 ;
        RECT 551.000000 269.850000 556.000000 270.150000 ;
        RECT 551.000000 285.850000 556.000000 286.150000 ;
        RECT 551.000000 301.850000 556.000000 302.150000 ;
        RECT 551.000000 297.850000 556.000000 298.150000 ;
        RECT 551.000000 293.850000 556.000000 294.150000 ;
        RECT 551.000000 289.850000 556.000000 290.150000 ;
        RECT 551.000000 309.850000 556.000000 310.150000 ;
        RECT 551.000000 313.850000 556.000000 314.150000 ;
        RECT 551.000000 317.850000 556.000000 318.150000 ;
        RECT 551.000000 321.850000 556.000000 322.150000 ;
        RECT 551.000000 325.850000 556.000000 326.150000 ;
        RECT 551.000000 329.850000 556.000000 330.150000 ;
        RECT 551.000000 333.850000 556.000000 334.150000 ;
        RECT 551.000000 337.850000 556.000000 338.150000 ;
        RECT 551.000000 341.850000 556.000000 342.150000 ;
        RECT 601.000000 1.850000 606.000000 2.150000 ;
        RECT 601.000000 5.850000 606.000000 6.150000 ;
        RECT 651.000000 1.850000 656.000000 2.150000 ;
        RECT 651.000000 5.850000 656.000000 6.150000 ;
        RECT 701.000000 1.850000 706.000000 2.150000 ;
        RECT 701.000000 5.850000 706.000000 6.150000 ;
        RECT 751.000000 1.850000 756.000000 2.150000 ;
        RECT 751.000000 5.850000 756.000000 6.150000 ;
        RECT 801.000000 1.850000 806.000000 2.150000 ;
        RECT 801.000000 5.850000 806.000000 6.150000 ;
        RECT 851.000000 1.850000 856.000000 2.150000 ;
        RECT 851.000000 5.850000 856.000000 6.150000 ;
        RECT 901.000000 1.850000 906.000000 2.150000 ;
        RECT 901.000000 5.850000 906.000000 6.150000 ;
        RECT 951.000000 1.850000 956.000000 2.150000 ;
        RECT 951.000000 5.850000 956.000000 6.150000 ;
        RECT 1001.000000 1.850000 1006.000000 2.150000 ;
        RECT 1001.000000 5.850000 1006.000000 6.150000 ;
        RECT 1051.000000 1.850000 1056.000000 2.150000 ;
        RECT 1051.000000 5.850000 1056.000000 6.150000 ;
        RECT 1101.000000 1.850000 1106.000000 2.150000 ;
        RECT 1101.000000 5.850000 1106.000000 6.150000 ;
        RECT 1151.000000 5.850000 1156.000000 6.150000 ;
        RECT 1172.000000 5.850000 1182.000000 6.150000 ;
        RECT 1151.000000 1.850000 1156.000000 2.150000 ;
        RECT 1172.000000 17.850000 1182.000000 18.150000 ;
        RECT 1172.000000 13.850000 1182.000000 14.150000 ;
        RECT 1172.000000 9.850000 1182.000000 10.150000 ;
        RECT 1172.000000 21.850000 1182.000000 22.150000 ;
        RECT 1172.000000 25.850000 1182.000000 26.150000 ;
        RECT 1172.000000 33.850000 1182.000000 34.150000 ;
        RECT 1172.000000 29.850000 1182.000000 30.150000 ;
        RECT 1172.000000 41.850000 1182.000000 42.150000 ;
        RECT 1172.000000 37.850000 1182.000000 38.150000 ;
        RECT 1172.000000 45.850000 1182.000000 46.150000 ;
        RECT 601.000000 261.850000 606.000000 262.150000 ;
        RECT 601.000000 265.850000 606.000000 266.150000 ;
        RECT 651.000000 261.850000 656.000000 262.150000 ;
        RECT 651.000000 265.850000 656.000000 266.150000 ;
        RECT 701.000000 265.850000 706.000000 266.150000 ;
        RECT 701.000000 261.850000 706.000000 262.150000 ;
        RECT 601.000000 305.850000 606.000000 306.150000 ;
        RECT 651.000000 305.850000 656.000000 306.150000 ;
        RECT 601.000000 277.850000 606.000000 278.150000 ;
        RECT 601.000000 269.850000 606.000000 270.150000 ;
        RECT 601.000000 273.850000 606.000000 274.150000 ;
        RECT 601.000000 281.850000 606.000000 282.150000 ;
        RECT 601.000000 285.850000 606.000000 286.150000 ;
        RECT 601.000000 289.850000 606.000000 290.150000 ;
        RECT 601.000000 293.850000 606.000000 294.150000 ;
        RECT 601.000000 297.850000 606.000000 298.150000 ;
        RECT 601.000000 301.850000 606.000000 302.150000 ;
        RECT 651.000000 277.850000 656.000000 278.150000 ;
        RECT 651.000000 273.850000 656.000000 274.150000 ;
        RECT 651.000000 269.850000 656.000000 270.150000 ;
        RECT 651.000000 281.850000 656.000000 282.150000 ;
        RECT 651.000000 285.850000 656.000000 286.150000 ;
        RECT 651.000000 289.850000 656.000000 290.150000 ;
        RECT 651.000000 293.850000 656.000000 294.150000 ;
        RECT 651.000000 301.850000 656.000000 302.150000 ;
        RECT 651.000000 297.850000 656.000000 298.150000 ;
        RECT 601.000000 321.850000 606.000000 322.150000 ;
        RECT 601.000000 317.850000 606.000000 318.150000 ;
        RECT 601.000000 309.850000 606.000000 310.150000 ;
        RECT 601.000000 313.850000 606.000000 314.150000 ;
        RECT 601.000000 325.850000 606.000000 326.150000 ;
        RECT 601.000000 329.850000 606.000000 330.150000 ;
        RECT 601.000000 333.850000 606.000000 334.150000 ;
        RECT 601.000000 337.850000 606.000000 338.150000 ;
        RECT 601.000000 341.850000 606.000000 342.150000 ;
        RECT 651.000000 313.850000 656.000000 314.150000 ;
        RECT 651.000000 309.850000 656.000000 310.150000 ;
        RECT 651.000000 321.850000 656.000000 322.150000 ;
        RECT 651.000000 317.850000 656.000000 318.150000 ;
        RECT 651.000000 329.850000 656.000000 330.150000 ;
        RECT 651.000000 325.850000 656.000000 326.150000 ;
        RECT 651.000000 333.850000 656.000000 334.150000 ;
        RECT 651.000000 337.850000 656.000000 338.150000 ;
        RECT 651.000000 341.850000 656.000000 342.150000 ;
        RECT 701.000000 305.850000 706.000000 306.150000 ;
        RECT 701.000000 281.850000 706.000000 282.150000 ;
        RECT 701.000000 277.850000 706.000000 278.150000 ;
        RECT 701.000000 273.850000 706.000000 274.150000 ;
        RECT 701.000000 269.850000 706.000000 270.150000 ;
        RECT 701.000000 285.850000 706.000000 286.150000 ;
        RECT 701.000000 301.850000 706.000000 302.150000 ;
        RECT 701.000000 297.850000 706.000000 298.150000 ;
        RECT 701.000000 293.850000 706.000000 294.150000 ;
        RECT 701.000000 289.850000 706.000000 290.150000 ;
        RECT 701.000000 309.850000 706.000000 310.150000 ;
        RECT 701.000000 313.850000 706.000000 314.150000 ;
        RECT 701.000000 317.850000 706.000000 318.150000 ;
        RECT 701.000000 321.850000 706.000000 322.150000 ;
        RECT 701.000000 325.850000 706.000000 326.150000 ;
        RECT 701.000000 329.850000 706.000000 330.150000 ;
        RECT 701.000000 333.850000 706.000000 334.150000 ;
        RECT 701.000000 337.850000 706.000000 338.150000 ;
        RECT 701.000000 341.850000 706.000000 342.150000 ;
        RECT 751.000000 261.850000 756.000000 262.150000 ;
        RECT 751.000000 265.850000 756.000000 266.150000 ;
        RECT 801.000000 261.850000 806.000000 262.150000 ;
        RECT 801.000000 265.850000 806.000000 266.150000 ;
        RECT 851.000000 265.850000 856.000000 266.150000 ;
        RECT 851.000000 261.850000 856.000000 262.150000 ;
        RECT 801.000000 305.850000 806.000000 306.150000 ;
        RECT 751.000000 305.850000 756.000000 306.150000 ;
        RECT 751.000000 285.850000 756.000000 286.150000 ;
        RECT 751.000000 281.850000 756.000000 282.150000 ;
        RECT 751.000000 269.850000 756.000000 270.150000 ;
        RECT 751.000000 273.850000 756.000000 274.150000 ;
        RECT 751.000000 277.850000 756.000000 278.150000 ;
        RECT 751.000000 289.850000 756.000000 290.150000 ;
        RECT 751.000000 293.850000 756.000000 294.150000 ;
        RECT 751.000000 297.850000 756.000000 298.150000 ;
        RECT 751.000000 301.850000 756.000000 302.150000 ;
        RECT 801.000000 277.850000 806.000000 278.150000 ;
        RECT 801.000000 269.850000 806.000000 270.150000 ;
        RECT 801.000000 273.850000 806.000000 274.150000 ;
        RECT 801.000000 281.850000 806.000000 282.150000 ;
        RECT 801.000000 285.850000 806.000000 286.150000 ;
        RECT 801.000000 289.850000 806.000000 290.150000 ;
        RECT 801.000000 293.850000 806.000000 294.150000 ;
        RECT 801.000000 301.850000 806.000000 302.150000 ;
        RECT 801.000000 297.850000 806.000000 298.150000 ;
        RECT 751.000000 321.850000 756.000000 322.150000 ;
        RECT 751.000000 317.850000 756.000000 318.150000 ;
        RECT 751.000000 309.850000 756.000000 310.150000 ;
        RECT 751.000000 313.850000 756.000000 314.150000 ;
        RECT 751.000000 325.850000 756.000000 326.150000 ;
        RECT 751.000000 329.850000 756.000000 330.150000 ;
        RECT 751.000000 333.850000 756.000000 334.150000 ;
        RECT 751.000000 337.850000 756.000000 338.150000 ;
        RECT 751.000000 341.850000 756.000000 342.150000 ;
        RECT 801.000000 313.850000 806.000000 314.150000 ;
        RECT 801.000000 309.850000 806.000000 310.150000 ;
        RECT 801.000000 321.850000 806.000000 322.150000 ;
        RECT 801.000000 317.850000 806.000000 318.150000 ;
        RECT 801.000000 329.850000 806.000000 330.150000 ;
        RECT 801.000000 325.850000 806.000000 326.150000 ;
        RECT 801.000000 333.850000 806.000000 334.150000 ;
        RECT 801.000000 337.850000 806.000000 338.150000 ;
        RECT 801.000000 341.850000 806.000000 342.150000 ;
        RECT 851.000000 305.850000 856.000000 306.150000 ;
        RECT 851.000000 281.850000 856.000000 282.150000 ;
        RECT 851.000000 277.850000 856.000000 278.150000 ;
        RECT 851.000000 273.850000 856.000000 274.150000 ;
        RECT 851.000000 269.850000 856.000000 270.150000 ;
        RECT 851.000000 285.850000 856.000000 286.150000 ;
        RECT 851.000000 301.850000 856.000000 302.150000 ;
        RECT 851.000000 297.850000 856.000000 298.150000 ;
        RECT 851.000000 293.850000 856.000000 294.150000 ;
        RECT 851.000000 289.850000 856.000000 290.150000 ;
        RECT 851.000000 309.850000 856.000000 310.150000 ;
        RECT 851.000000 313.850000 856.000000 314.150000 ;
        RECT 851.000000 317.850000 856.000000 318.150000 ;
        RECT 851.000000 321.850000 856.000000 322.150000 ;
        RECT 851.000000 325.850000 856.000000 326.150000 ;
        RECT 851.000000 329.850000 856.000000 330.150000 ;
        RECT 851.000000 333.850000 856.000000 334.150000 ;
        RECT 851.000000 337.850000 856.000000 338.150000 ;
        RECT 851.000000 341.850000 856.000000 342.150000 ;
        RECT 1172.000000 61.850000 1182.000000 62.150000 ;
        RECT 1172.000000 57.850000 1182.000000 58.150000 ;
        RECT 1172.000000 53.850000 1182.000000 54.150000 ;
        RECT 1172.000000 49.850000 1182.000000 50.150000 ;
        RECT 1172.000000 73.850000 1182.000000 74.150000 ;
        RECT 1172.000000 69.850000 1182.000000 70.150000 ;
        RECT 1172.000000 65.850000 1182.000000 66.150000 ;
        RECT 1172.000000 77.850000 1182.000000 78.150000 ;
        RECT 1172.000000 81.850000 1182.000000 82.150000 ;
        RECT 1172.000000 101.850000 1182.000000 102.150000 ;
        RECT 1172.000000 89.850000 1182.000000 90.150000 ;
        RECT 1172.000000 85.850000 1182.000000 86.150000 ;
        RECT 1172.000000 93.850000 1182.000000 94.150000 ;
        RECT 1172.000000 97.850000 1182.000000 98.150000 ;
        RECT 1172.000000 117.850000 1182.000000 118.150000 ;
        RECT 1172.000000 113.850000 1182.000000 114.150000 ;
        RECT 1172.000000 105.850000 1182.000000 106.150000 ;
        RECT 1172.000000 109.850000 1182.000000 110.150000 ;
        RECT 1151.000000 133.850000 1156.000000 134.150000 ;
        RECT 1172.000000 129.850000 1182.000000 130.150000 ;
        RECT 1172.000000 125.850000 1182.000000 126.150000 ;
        RECT 1172.000000 121.850000 1182.000000 122.150000 ;
        RECT 1172.000000 133.850000 1182.000000 134.150000 ;
        RECT 1172.000000 137.850000 1182.000000 138.150000 ;
        RECT 1172.000000 141.850000 1182.000000 142.150000 ;
        RECT 1172.000000 145.850000 1182.000000 146.150000 ;
        RECT 1172.000000 149.850000 1182.000000 150.150000 ;
        RECT 1172.000000 153.850000 1182.000000 154.150000 ;
        RECT 1172.000000 165.850000 1182.000000 166.150000 ;
        RECT 1172.000000 161.850000 1182.000000 162.150000 ;
        RECT 1172.000000 157.850000 1182.000000 158.150000 ;
        RECT 1172.000000 169.850000 1182.000000 170.150000 ;
        RECT 1172.000000 173.850000 1182.000000 174.150000 ;
        RECT 1172.000000 177.850000 1182.000000 178.150000 ;
        RECT 1172.000000 181.850000 1182.000000 182.150000 ;
        RECT 1172.000000 185.850000 1182.000000 186.150000 ;
        RECT 1172.000000 189.850000 1182.000000 190.150000 ;
        RECT 1172.000000 193.850000 1182.000000 194.150000 ;
        RECT 901.000000 261.850000 906.000000 262.150000 ;
        RECT 901.000000 265.850000 906.000000 266.150000 ;
        RECT 951.000000 265.850000 956.000000 266.150000 ;
        RECT 951.000000 261.850000 956.000000 262.150000 ;
        RECT 1001.000000 261.850000 1006.000000 262.150000 ;
        RECT 1001.000000 265.850000 1006.000000 266.150000 ;
        RECT 951.000000 305.850000 956.000000 306.150000 ;
        RECT 901.000000 305.850000 906.000000 306.150000 ;
        RECT 901.000000 285.850000 906.000000 286.150000 ;
        RECT 901.000000 281.850000 906.000000 282.150000 ;
        RECT 901.000000 269.850000 906.000000 270.150000 ;
        RECT 901.000000 273.850000 906.000000 274.150000 ;
        RECT 901.000000 277.850000 906.000000 278.150000 ;
        RECT 901.000000 289.850000 906.000000 290.150000 ;
        RECT 901.000000 293.850000 906.000000 294.150000 ;
        RECT 901.000000 297.850000 906.000000 298.150000 ;
        RECT 901.000000 301.850000 906.000000 302.150000 ;
        RECT 951.000000 269.850000 956.000000 270.150000 ;
        RECT 951.000000 273.850000 956.000000 274.150000 ;
        RECT 951.000000 277.850000 956.000000 278.150000 ;
        RECT 951.000000 281.850000 956.000000 282.150000 ;
        RECT 951.000000 285.850000 956.000000 286.150000 ;
        RECT 951.000000 301.850000 956.000000 302.150000 ;
        RECT 951.000000 297.850000 956.000000 298.150000 ;
        RECT 951.000000 293.850000 956.000000 294.150000 ;
        RECT 951.000000 289.850000 956.000000 290.150000 ;
        RECT 901.000000 321.850000 906.000000 322.150000 ;
        RECT 901.000000 309.850000 906.000000 310.150000 ;
        RECT 901.000000 313.850000 906.000000 314.150000 ;
        RECT 901.000000 317.850000 906.000000 318.150000 ;
        RECT 901.000000 325.850000 906.000000 326.150000 ;
        RECT 901.000000 329.850000 906.000000 330.150000 ;
        RECT 901.000000 333.850000 906.000000 334.150000 ;
        RECT 901.000000 337.850000 906.000000 338.150000 ;
        RECT 901.000000 341.850000 906.000000 342.150000 ;
        RECT 951.000000 313.850000 956.000000 314.150000 ;
        RECT 951.000000 309.850000 956.000000 310.150000 ;
        RECT 951.000000 317.850000 956.000000 318.150000 ;
        RECT 951.000000 321.850000 956.000000 322.150000 ;
        RECT 951.000000 325.850000 956.000000 326.150000 ;
        RECT 951.000000 329.850000 956.000000 330.150000 ;
        RECT 951.000000 333.850000 956.000000 334.150000 ;
        RECT 951.000000 337.850000 956.000000 338.150000 ;
        RECT 951.000000 341.850000 956.000000 342.150000 ;
        RECT 1001.000000 305.850000 1006.000000 306.150000 ;
        RECT 1001.000000 277.850000 1006.000000 278.150000 ;
        RECT 1001.000000 269.850000 1006.000000 270.150000 ;
        RECT 1001.000000 273.850000 1006.000000 274.150000 ;
        RECT 1001.000000 285.850000 1006.000000 286.150000 ;
        RECT 1001.000000 281.850000 1006.000000 282.150000 ;
        RECT 1001.000000 289.850000 1006.000000 290.150000 ;
        RECT 1001.000000 293.850000 1006.000000 294.150000 ;
        RECT 1001.000000 301.850000 1006.000000 302.150000 ;
        RECT 1001.000000 297.850000 1006.000000 298.150000 ;
        RECT 1001.000000 313.850000 1006.000000 314.150000 ;
        RECT 1001.000000 309.850000 1006.000000 310.150000 ;
        RECT 1001.000000 317.850000 1006.000000 318.150000 ;
        RECT 1001.000000 321.850000 1006.000000 322.150000 ;
        RECT 1001.000000 329.850000 1006.000000 330.150000 ;
        RECT 1001.000000 325.850000 1006.000000 326.150000 ;
        RECT 1001.000000 333.850000 1006.000000 334.150000 ;
        RECT 1001.000000 337.850000 1006.000000 338.150000 ;
        RECT 1001.000000 341.850000 1006.000000 342.150000 ;
        RECT 1051.000000 261.850000 1056.000000 262.150000 ;
        RECT 1051.000000 265.850000 1056.000000 266.150000 ;
        RECT 1101.000000 265.850000 1106.000000 266.150000 ;
        RECT 1101.000000 261.850000 1106.000000 262.150000 ;
        RECT 1172.000000 197.850000 1182.000000 198.150000 ;
        RECT 1172.000000 201.850000 1182.000000 202.150000 ;
        RECT 1172.000000 205.850000 1182.000000 206.150000 ;
        RECT 1172.000000 209.850000 1182.000000 210.150000 ;
        RECT 1172.000000 221.850000 1182.000000 222.150000 ;
        RECT 1172.000000 217.850000 1182.000000 218.150000 ;
        RECT 1172.000000 213.850000 1182.000000 214.150000 ;
        RECT 1172.000000 225.850000 1182.000000 226.150000 ;
        RECT 1172.000000 229.850000 1182.000000 230.150000 ;
        RECT 1172.000000 233.850000 1182.000000 234.150000 ;
        RECT 1172.000000 237.850000 1182.000000 238.150000 ;
        RECT 1172.000000 241.850000 1182.000000 242.150000 ;
        RECT 1172.000000 245.850000 1182.000000 246.150000 ;
        RECT 1172.000000 249.850000 1182.000000 250.150000 ;
        RECT 1151.000000 257.850000 1156.000000 258.150000 ;
        RECT 1151.000000 265.850000 1156.000000 266.150000 ;
        RECT 1151.000000 261.850000 1156.000000 262.150000 ;
        RECT 1172.000000 265.850000 1182.000000 266.150000 ;
        RECT 1172.000000 253.850000 1182.000000 254.150000 ;
        RECT 1172.000000 257.850000 1182.000000 258.150000 ;
        RECT 1172.000000 261.850000 1182.000000 262.150000 ;
        RECT 1101.000000 305.850000 1106.000000 306.150000 ;
        RECT 1051.000000 305.850000 1056.000000 306.150000 ;
        RECT 1051.000000 285.850000 1056.000000 286.150000 ;
        RECT 1051.000000 281.850000 1056.000000 282.150000 ;
        RECT 1051.000000 273.850000 1056.000000 274.150000 ;
        RECT 1051.000000 269.850000 1056.000000 270.150000 ;
        RECT 1051.000000 277.850000 1056.000000 278.150000 ;
        RECT 1051.000000 289.850000 1056.000000 290.150000 ;
        RECT 1051.000000 293.850000 1056.000000 294.150000 ;
        RECT 1051.000000 297.850000 1056.000000 298.150000 ;
        RECT 1051.000000 301.850000 1056.000000 302.150000 ;
        RECT 1101.000000 269.850000 1106.000000 270.150000 ;
        RECT 1101.000000 273.850000 1106.000000 274.150000 ;
        RECT 1101.000000 277.850000 1106.000000 278.150000 ;
        RECT 1101.000000 281.850000 1106.000000 282.150000 ;
        RECT 1101.000000 285.850000 1106.000000 286.150000 ;
        RECT 1101.000000 301.850000 1106.000000 302.150000 ;
        RECT 1101.000000 297.850000 1106.000000 298.150000 ;
        RECT 1101.000000 293.850000 1106.000000 294.150000 ;
        RECT 1101.000000 289.850000 1106.000000 290.150000 ;
        RECT 1051.000000 321.850000 1056.000000 322.150000 ;
        RECT 1051.000000 309.850000 1056.000000 310.150000 ;
        RECT 1051.000000 313.850000 1056.000000 314.150000 ;
        RECT 1051.000000 317.850000 1056.000000 318.150000 ;
        RECT 1051.000000 325.850000 1056.000000 326.150000 ;
        RECT 1051.000000 329.850000 1056.000000 330.150000 ;
        RECT 1051.000000 333.850000 1056.000000 334.150000 ;
        RECT 1051.000000 337.850000 1056.000000 338.150000 ;
        RECT 1051.000000 341.850000 1056.000000 342.150000 ;
        RECT 1101.000000 313.850000 1106.000000 314.150000 ;
        RECT 1101.000000 309.850000 1106.000000 310.150000 ;
        RECT 1101.000000 317.850000 1106.000000 318.150000 ;
        RECT 1101.000000 321.850000 1106.000000 322.150000 ;
        RECT 1101.000000 325.850000 1106.000000 326.150000 ;
        RECT 1101.000000 329.850000 1106.000000 330.150000 ;
        RECT 1101.000000 333.850000 1106.000000 334.150000 ;
        RECT 1101.000000 337.850000 1106.000000 338.150000 ;
        RECT 1101.000000 341.850000 1106.000000 342.150000 ;
        RECT 1151.000000 305.850000 1156.000000 306.150000 ;
        RECT 1172.000000 305.850000 1182.000000 306.150000 ;
        RECT 1151.000000 277.850000 1156.000000 278.150000 ;
        RECT 1151.000000 269.850000 1156.000000 270.150000 ;
        RECT 1151.000000 273.850000 1156.000000 274.150000 ;
        RECT 1151.000000 281.850000 1156.000000 282.150000 ;
        RECT 1151.000000 285.850000 1156.000000 286.150000 ;
        RECT 1172.000000 277.850000 1182.000000 278.150000 ;
        RECT 1172.000000 269.850000 1182.000000 270.150000 ;
        RECT 1172.000000 273.850000 1182.000000 274.150000 ;
        RECT 1172.000000 281.850000 1182.000000 282.150000 ;
        RECT 1172.000000 285.850000 1182.000000 286.150000 ;
        RECT 1151.000000 301.850000 1156.000000 302.150000 ;
        RECT 1151.000000 297.850000 1156.000000 298.150000 ;
        RECT 1151.000000 289.850000 1156.000000 290.150000 ;
        RECT 1151.000000 293.850000 1156.000000 294.150000 ;
        RECT 1172.000000 301.850000 1182.000000 302.150000 ;
        RECT 1172.000000 289.850000 1182.000000 290.150000 ;
        RECT 1172.000000 293.850000 1182.000000 294.150000 ;
        RECT 1172.000000 297.850000 1182.000000 298.150000 ;
        RECT 1151.000000 321.850000 1156.000000 322.150000 ;
        RECT 1151.000000 317.850000 1156.000000 318.150000 ;
        RECT 1151.000000 309.850000 1156.000000 310.150000 ;
        RECT 1151.000000 313.850000 1156.000000 314.150000 ;
        RECT 1172.000000 321.850000 1182.000000 322.150000 ;
        RECT 1172.000000 309.850000 1182.000000 310.150000 ;
        RECT 1172.000000 313.850000 1182.000000 314.150000 ;
        RECT 1172.000000 317.850000 1182.000000 318.150000 ;
        RECT 1151.000000 329.850000 1156.000000 330.150000 ;
        RECT 1151.000000 325.850000 1156.000000 326.150000 ;
        RECT 1151.000000 333.850000 1156.000000 334.150000 ;
        RECT 1151.000000 337.850000 1156.000000 338.150000 ;
        RECT 1151.000000 341.850000 1156.000000 342.150000 ;
        RECT 1172.000000 329.850000 1182.000000 330.150000 ;
        RECT 1172.000000 325.850000 1182.000000 326.150000 ;
        RECT 1172.000000 333.850000 1182.000000 334.150000 ;
        RECT 1172.000000 337.850000 1182.000000 338.150000 ;
        RECT 1172.000000 341.850000 1182.000000 342.150000 ;
        RECT 4.000000 357.850000 14.000000 358.150000 ;
        RECT 4.000000 353.850000 14.000000 354.150000 ;
        RECT 4.000000 345.850000 14.000000 346.150000 ;
        RECT 4.000000 349.850000 14.000000 350.150000 ;
        RECT 4.000000 369.850000 14.000000 370.150000 ;
        RECT 4.000000 365.850000 14.000000 366.150000 ;
        RECT 4.000000 361.850000 14.000000 362.150000 ;
        RECT 4.000000 377.850000 14.000000 378.150000 ;
        RECT 4.000000 373.850000 14.000000 374.150000 ;
        RECT 51.000000 345.850000 56.000000 346.150000 ;
        RECT 51.000000 369.850000 56.000000 370.150000 ;
        RECT 51.000000 365.850000 56.000000 366.150000 ;
        RECT 51.000000 361.850000 56.000000 362.150000 ;
        RECT 51.000000 373.850000 56.000000 374.150000 ;
        RECT 51.000000 377.850000 56.000000 378.150000 ;
        RECT 4.000000 393.850000 14.000000 394.150000 ;
        RECT 4.000000 389.850000 14.000000 390.150000 ;
        RECT 4.000000 381.850000 14.000000 382.150000 ;
        RECT 4.000000 385.850000 14.000000 386.150000 ;
        RECT 4.000000 397.850000 14.000000 398.150000 ;
        RECT 4.000000 401.850000 14.000000 402.150000 ;
        RECT 4.000000 405.850000 14.000000 406.150000 ;
        RECT 4.000000 409.850000 14.000000 410.150000 ;
        RECT 4.000000 413.850000 14.000000 414.150000 ;
        RECT 51.000000 397.850000 56.000000 398.150000 ;
        RECT 51.000000 385.850000 56.000000 386.150000 ;
        RECT 51.000000 381.850000 56.000000 382.150000 ;
        RECT 51.000000 389.850000 56.000000 390.150000 ;
        RECT 51.000000 393.850000 56.000000 394.150000 ;
        RECT 51.000000 413.850000 56.000000 414.150000 ;
        RECT 51.000000 409.850000 56.000000 410.150000 ;
        RECT 51.000000 405.850000 56.000000 406.150000 ;
        RECT 51.000000 401.850000 56.000000 402.150000 ;
        RECT 101.000000 345.850000 106.000000 346.150000 ;
        RECT 101.000000 349.850000 106.000000 350.150000 ;
        RECT 101.000000 353.850000 106.000000 354.150000 ;
        RECT 101.000000 357.850000 106.000000 358.150000 ;
        RECT 101.000000 361.850000 106.000000 362.150000 ;
        RECT 101.000000 365.850000 106.000000 366.150000 ;
        RECT 101.000000 369.850000 106.000000 370.150000 ;
        RECT 101.000000 373.850000 106.000000 374.150000 ;
        RECT 101.000000 377.850000 106.000000 378.150000 ;
        RECT 101.000000 397.850000 106.000000 398.150000 ;
        RECT 101.000000 381.850000 106.000000 382.150000 ;
        RECT 101.000000 385.850000 106.000000 386.150000 ;
        RECT 101.000000 389.850000 106.000000 390.150000 ;
        RECT 101.000000 393.850000 106.000000 394.150000 ;
        RECT 101.000000 413.850000 106.000000 414.150000 ;
        RECT 101.000000 409.850000 106.000000 410.150000 ;
        RECT 101.000000 405.850000 106.000000 406.150000 ;
        RECT 101.000000 401.850000 106.000000 402.150000 ;
        RECT 4.000000 433.850000 14.000000 434.150000 ;
        RECT 4.000000 429.850000 14.000000 430.150000 ;
        RECT 4.000000 421.850000 14.000000 422.150000 ;
        RECT 4.000000 417.850000 14.000000 418.150000 ;
        RECT 4.000000 425.850000 14.000000 426.150000 ;
        RECT 4.000000 437.850000 14.000000 438.150000 ;
        RECT 4.000000 441.850000 14.000000 442.150000 ;
        RECT 4.000000 445.850000 14.000000 446.150000 ;
        RECT 4.000000 449.850000 14.000000 450.150000 ;
        RECT 4.000000 453.850000 14.000000 454.150000 ;
        RECT 51.000000 417.850000 56.000000 418.150000 ;
        RECT 51.000000 421.850000 56.000000 422.150000 ;
        RECT 51.000000 425.850000 56.000000 426.150000 ;
        RECT 51.000000 429.850000 56.000000 430.150000 ;
        RECT 51.000000 433.850000 56.000000 434.150000 ;
        RECT 51.000000 453.850000 56.000000 454.150000 ;
        RECT 51.000000 449.850000 56.000000 450.150000 ;
        RECT 51.000000 445.850000 56.000000 446.150000 ;
        RECT 51.000000 441.850000 56.000000 442.150000 ;
        RECT 51.000000 437.850000 56.000000 438.150000 ;
        RECT 4.000000 469.850000 14.000000 470.150000 ;
        RECT 4.000000 465.850000 14.000000 466.150000 ;
        RECT 4.000000 457.850000 14.000000 458.150000 ;
        RECT 4.000000 461.850000 14.000000 462.150000 ;
        RECT 4.000000 473.850000 14.000000 474.150000 ;
        RECT 4.000000 477.850000 14.000000 478.150000 ;
        RECT 4.000000 481.850000 14.000000 482.150000 ;
        RECT 4.000000 485.850000 14.000000 486.150000 ;
        RECT 4.000000 489.850000 14.000000 490.150000 ;
        RECT 51.000000 461.850000 56.000000 462.150000 ;
        RECT 51.000000 457.850000 56.000000 458.150000 ;
        RECT 51.000000 465.850000 56.000000 466.150000 ;
        RECT 51.000000 469.850000 56.000000 470.150000 ;
        RECT 51.000000 489.850000 56.000000 490.150000 ;
        RECT 51.000000 485.850000 56.000000 486.150000 ;
        RECT 51.000000 481.850000 56.000000 482.150000 ;
        RECT 51.000000 477.850000 56.000000 478.150000 ;
        RECT 51.000000 473.850000 56.000000 474.150000 ;
        RECT 101.000000 433.850000 106.000000 434.150000 ;
        RECT 101.000000 417.850000 106.000000 418.150000 ;
        RECT 101.000000 421.850000 106.000000 422.150000 ;
        RECT 101.000000 425.850000 106.000000 426.150000 ;
        RECT 101.000000 429.850000 106.000000 430.150000 ;
        RECT 101.000000 437.850000 106.000000 438.150000 ;
        RECT 101.000000 441.850000 106.000000 442.150000 ;
        RECT 101.000000 445.850000 106.000000 446.150000 ;
        RECT 101.000000 449.850000 106.000000 450.150000 ;
        RECT 101.000000 453.850000 106.000000 454.150000 ;
        RECT 101.000000 469.850000 106.000000 470.150000 ;
        RECT 101.000000 465.850000 106.000000 466.150000 ;
        RECT 101.000000 461.850000 106.000000 462.150000 ;
        RECT 101.000000 457.850000 106.000000 458.150000 ;
        RECT 101.000000 473.850000 106.000000 474.150000 ;
        RECT 101.000000 477.850000 106.000000 478.150000 ;
        RECT 101.000000 481.850000 106.000000 482.150000 ;
        RECT 101.000000 485.850000 106.000000 486.150000 ;
        RECT 101.000000 489.850000 106.000000 490.150000 ;
        RECT 151.000000 349.850000 156.000000 350.150000 ;
        RECT 151.000000 345.850000 156.000000 346.150000 ;
        RECT 151.000000 353.850000 156.000000 354.150000 ;
        RECT 151.000000 357.850000 156.000000 358.150000 ;
        RECT 151.000000 361.850000 156.000000 362.150000 ;
        RECT 151.000000 365.850000 156.000000 366.150000 ;
        RECT 151.000000 369.850000 156.000000 370.150000 ;
        RECT 151.000000 373.850000 156.000000 374.150000 ;
        RECT 151.000000 377.850000 156.000000 378.150000 ;
        RECT 201.000000 349.850000 206.000000 350.150000 ;
        RECT 201.000000 345.850000 206.000000 346.150000 ;
        RECT 201.000000 353.850000 206.000000 354.150000 ;
        RECT 201.000000 357.850000 206.000000 358.150000 ;
        RECT 201.000000 377.850000 206.000000 378.150000 ;
        RECT 201.000000 373.850000 206.000000 374.150000 ;
        RECT 201.000000 369.850000 206.000000 370.150000 ;
        RECT 201.000000 365.850000 206.000000 366.150000 ;
        RECT 201.000000 361.850000 206.000000 362.150000 ;
        RECT 151.000000 385.850000 156.000000 386.150000 ;
        RECT 151.000000 381.850000 156.000000 382.150000 ;
        RECT 151.000000 393.850000 156.000000 394.150000 ;
        RECT 151.000000 389.850000 156.000000 390.150000 ;
        RECT 151.000000 397.850000 156.000000 398.150000 ;
        RECT 151.000000 401.850000 156.000000 402.150000 ;
        RECT 201.000000 381.850000 206.000000 382.150000 ;
        RECT 201.000000 385.850000 206.000000 386.150000 ;
        RECT 201.000000 397.850000 206.000000 398.150000 ;
        RECT 201.000000 393.850000 206.000000 394.150000 ;
        RECT 201.000000 389.850000 206.000000 390.150000 ;
        RECT 201.000000 413.850000 206.000000 414.150000 ;
        RECT 201.000000 409.850000 206.000000 410.150000 ;
        RECT 201.000000 405.850000 206.000000 406.150000 ;
        RECT 201.000000 401.850000 206.000000 402.150000 ;
        RECT 251.000000 345.850000 256.000000 346.150000 ;
        RECT 251.000000 349.850000 256.000000 350.150000 ;
        RECT 251.000000 353.850000 256.000000 354.150000 ;
        RECT 251.000000 357.850000 256.000000 358.150000 ;
        RECT 251.000000 365.850000 256.000000 366.150000 ;
        RECT 251.000000 361.850000 256.000000 362.150000 ;
        RECT 251.000000 369.850000 256.000000 370.150000 ;
        RECT 251.000000 373.850000 256.000000 374.150000 ;
        RECT 251.000000 377.850000 256.000000 378.150000 ;
        RECT 251.000000 381.850000 256.000000 382.150000 ;
        RECT 251.000000 385.850000 256.000000 386.150000 ;
        RECT 251.000000 393.850000 256.000000 394.150000 ;
        RECT 251.000000 389.850000 256.000000 390.150000 ;
        RECT 251.000000 397.850000 256.000000 398.150000 ;
        RECT 251.000000 401.850000 256.000000 402.150000 ;
        RECT 151.000000 453.850000 156.000000 454.150000 ;
        RECT 201.000000 429.850000 206.000000 430.150000 ;
        RECT 201.000000 425.850000 206.000000 426.150000 ;
        RECT 201.000000 421.850000 206.000000 422.150000 ;
        RECT 201.000000 417.850000 206.000000 418.150000 ;
        RECT 201.000000 433.850000 206.000000 434.150000 ;
        RECT 201.000000 453.850000 206.000000 454.150000 ;
        RECT 201.000000 449.850000 206.000000 450.150000 ;
        RECT 201.000000 445.850000 206.000000 446.150000 ;
        RECT 201.000000 441.850000 206.000000 442.150000 ;
        RECT 201.000000 437.850000 206.000000 438.150000 ;
        RECT 151.000000 461.850000 156.000000 462.150000 ;
        RECT 151.000000 457.850000 156.000000 458.150000 ;
        RECT 151.000000 469.850000 156.000000 470.150000 ;
        RECT 151.000000 465.850000 156.000000 466.150000 ;
        RECT 151.000000 481.850000 156.000000 482.150000 ;
        RECT 151.000000 477.850000 156.000000 478.150000 ;
        RECT 151.000000 473.850000 156.000000 474.150000 ;
        RECT 151.000000 489.850000 156.000000 490.150000 ;
        RECT 151.000000 485.850000 156.000000 486.150000 ;
        RECT 201.000000 461.850000 206.000000 462.150000 ;
        RECT 201.000000 457.850000 206.000000 458.150000 ;
        RECT 201.000000 465.850000 206.000000 466.150000 ;
        RECT 201.000000 469.850000 206.000000 470.150000 ;
        RECT 201.000000 489.850000 206.000000 490.150000 ;
        RECT 201.000000 485.850000 206.000000 486.150000 ;
        RECT 201.000000 481.850000 206.000000 482.150000 ;
        RECT 201.000000 477.850000 206.000000 478.150000 ;
        RECT 201.000000 473.850000 206.000000 474.150000 ;
        RECT 251.000000 453.850000 256.000000 454.150000 ;
        RECT 251.000000 457.850000 256.000000 458.150000 ;
        RECT 251.000000 461.850000 256.000000 462.150000 ;
        RECT 251.000000 465.850000 256.000000 466.150000 ;
        RECT 251.000000 469.850000 256.000000 470.150000 ;
        RECT 251.000000 481.850000 256.000000 482.150000 ;
        RECT 251.000000 473.850000 256.000000 474.150000 ;
        RECT 251.000000 477.850000 256.000000 478.150000 ;
        RECT 251.000000 485.850000 256.000000 486.150000 ;
        RECT 251.000000 489.850000 256.000000 490.150000 ;
        RECT 4.000000 505.850000 14.000000 506.150000 ;
        RECT 4.000000 501.850000 14.000000 502.150000 ;
        RECT 4.000000 497.850000 14.000000 498.150000 ;
        RECT 4.000000 493.850000 14.000000 494.150000 ;
        RECT 4.000000 513.850000 14.000000 514.150000 ;
        RECT 4.000000 509.850000 14.000000 510.150000 ;
        RECT 51.000000 493.850000 56.000000 494.150000 ;
        RECT 51.000000 497.850000 56.000000 498.150000 ;
        RECT 51.000000 501.850000 56.000000 502.150000 ;
        RECT 51.000000 505.850000 56.000000 506.150000 ;
        RECT 51.000000 513.850000 56.000000 514.150000 ;
        RECT 51.000000 509.850000 56.000000 510.150000 ;
        RECT 101.000000 505.850000 106.000000 506.150000 ;
        RECT 101.000000 501.850000 106.000000 502.150000 ;
        RECT 101.000000 497.850000 106.000000 498.150000 ;
        RECT 101.000000 493.850000 106.000000 494.150000 ;
        RECT 101.000000 513.850000 106.000000 514.150000 ;
        RECT 101.000000 509.850000 106.000000 510.150000 ;
        RECT 151.000000 493.850000 156.000000 494.150000 ;
        RECT 151.000000 497.850000 156.000000 498.150000 ;
        RECT 151.000000 501.850000 156.000000 502.150000 ;
        RECT 151.000000 505.850000 156.000000 506.150000 ;
        RECT 151.000000 513.850000 156.000000 514.150000 ;
        RECT 151.000000 509.850000 156.000000 510.150000 ;
        RECT 201.000000 497.850000 206.000000 498.150000 ;
        RECT 201.000000 493.850000 206.000000 494.150000 ;
        RECT 201.000000 501.850000 206.000000 502.150000 ;
        RECT 201.000000 505.850000 206.000000 506.150000 ;
        RECT 201.000000 513.850000 206.000000 514.150000 ;
        RECT 201.000000 509.850000 206.000000 510.150000 ;
        RECT 251.000000 493.850000 256.000000 494.150000 ;
        RECT 251.000000 497.850000 256.000000 498.150000 ;
        RECT 251.000000 501.850000 256.000000 502.150000 ;
        RECT 251.000000 505.850000 256.000000 506.150000 ;
        RECT 251.000000 513.850000 256.000000 514.150000 ;
        RECT 251.000000 509.850000 256.000000 510.150000 ;
        RECT 301.000000 345.850000 306.000000 346.150000 ;
        RECT 301.000000 349.850000 306.000000 350.150000 ;
        RECT 301.000000 353.850000 306.000000 354.150000 ;
        RECT 301.000000 357.850000 306.000000 358.150000 ;
        RECT 301.000000 369.850000 306.000000 370.150000 ;
        RECT 301.000000 365.850000 306.000000 366.150000 ;
        RECT 301.000000 361.850000 306.000000 362.150000 ;
        RECT 301.000000 377.850000 306.000000 378.150000 ;
        RECT 301.000000 373.850000 306.000000 374.150000 ;
        RECT 351.000000 349.850000 356.000000 350.150000 ;
        RECT 351.000000 345.850000 356.000000 346.150000 ;
        RECT 351.000000 353.850000 356.000000 354.150000 ;
        RECT 351.000000 357.850000 356.000000 358.150000 ;
        RECT 351.000000 377.850000 356.000000 378.150000 ;
        RECT 351.000000 373.850000 356.000000 374.150000 ;
        RECT 351.000000 369.850000 356.000000 370.150000 ;
        RECT 351.000000 365.850000 356.000000 366.150000 ;
        RECT 351.000000 361.850000 356.000000 362.150000 ;
        RECT 301.000000 385.850000 306.000000 386.150000 ;
        RECT 301.000000 381.850000 306.000000 382.150000 ;
        RECT 301.000000 397.850000 306.000000 398.150000 ;
        RECT 301.000000 389.850000 306.000000 390.150000 ;
        RECT 301.000000 393.850000 306.000000 394.150000 ;
        RECT 301.000000 405.850000 306.000000 406.150000 ;
        RECT 301.000000 401.850000 306.000000 402.150000 ;
        RECT 301.000000 413.850000 306.000000 414.150000 ;
        RECT 301.000000 409.850000 306.000000 410.150000 ;
        RECT 351.000000 381.850000 356.000000 382.150000 ;
        RECT 351.000000 385.850000 356.000000 386.150000 ;
        RECT 351.000000 393.850000 356.000000 394.150000 ;
        RECT 351.000000 389.850000 356.000000 390.150000 ;
        RECT 351.000000 397.850000 356.000000 398.150000 ;
        RECT 351.000000 413.850000 356.000000 414.150000 ;
        RECT 351.000000 409.850000 356.000000 410.150000 ;
        RECT 351.000000 405.850000 356.000000 406.150000 ;
        RECT 351.000000 401.850000 356.000000 402.150000 ;
        RECT 401.000000 357.850000 406.000000 358.150000 ;
        RECT 401.000000 353.850000 406.000000 354.150000 ;
        RECT 401.000000 349.850000 406.000000 350.150000 ;
        RECT 401.000000 345.850000 406.000000 346.150000 ;
        RECT 401.000000 361.850000 406.000000 362.150000 ;
        RECT 401.000000 365.850000 406.000000 366.150000 ;
        RECT 401.000000 369.850000 406.000000 370.150000 ;
        RECT 401.000000 377.850000 406.000000 378.150000 ;
        RECT 401.000000 373.850000 406.000000 374.150000 ;
        RECT 401.000000 385.850000 406.000000 386.150000 ;
        RECT 401.000000 381.850000 406.000000 382.150000 ;
        RECT 401.000000 393.850000 406.000000 394.150000 ;
        RECT 401.000000 389.850000 406.000000 390.150000 ;
        RECT 401.000000 397.850000 406.000000 398.150000 ;
        RECT 401.000000 401.850000 406.000000 402.150000 ;
        RECT 401.000000 405.850000 406.000000 406.150000 ;
        RECT 401.000000 409.850000 406.000000 410.150000 ;
        RECT 401.000000 413.850000 406.000000 414.150000 ;
        RECT 301.000000 425.850000 306.000000 426.150000 ;
        RECT 301.000000 417.850000 306.000000 418.150000 ;
        RECT 301.000000 421.850000 306.000000 422.150000 ;
        RECT 301.000000 429.850000 306.000000 430.150000 ;
        RECT 301.000000 433.850000 306.000000 434.150000 ;
        RECT 301.000000 441.850000 306.000000 442.150000 ;
        RECT 301.000000 437.850000 306.000000 438.150000 ;
        RECT 301.000000 453.850000 306.000000 454.150000 ;
        RECT 301.000000 449.850000 306.000000 450.150000 ;
        RECT 301.000000 445.850000 306.000000 446.150000 ;
        RECT 351.000000 417.850000 356.000000 418.150000 ;
        RECT 351.000000 421.850000 356.000000 422.150000 ;
        RECT 351.000000 425.850000 356.000000 426.150000 ;
        RECT 351.000000 429.850000 356.000000 430.150000 ;
        RECT 351.000000 433.850000 356.000000 434.150000 ;
        RECT 351.000000 437.850000 356.000000 438.150000 ;
        RECT 351.000000 441.850000 356.000000 442.150000 ;
        RECT 351.000000 445.850000 356.000000 446.150000 ;
        RECT 351.000000 449.850000 356.000000 450.150000 ;
        RECT 351.000000 453.850000 356.000000 454.150000 ;
        RECT 301.000000 461.850000 306.000000 462.150000 ;
        RECT 301.000000 457.850000 306.000000 458.150000 ;
        RECT 301.000000 465.850000 306.000000 466.150000 ;
        RECT 301.000000 469.850000 306.000000 470.150000 ;
        RECT 301.000000 481.850000 306.000000 482.150000 ;
        RECT 301.000000 477.850000 306.000000 478.150000 ;
        RECT 301.000000 473.850000 306.000000 474.150000 ;
        RECT 301.000000 489.850000 306.000000 490.150000 ;
        RECT 301.000000 485.850000 306.000000 486.150000 ;
        RECT 351.000000 461.850000 356.000000 462.150000 ;
        RECT 351.000000 457.850000 356.000000 458.150000 ;
        RECT 351.000000 465.850000 356.000000 466.150000 ;
        RECT 351.000000 469.850000 356.000000 470.150000 ;
        RECT 351.000000 481.850000 356.000000 482.150000 ;
        RECT 351.000000 473.850000 356.000000 474.150000 ;
        RECT 351.000000 477.850000 356.000000 478.150000 ;
        RECT 351.000000 485.850000 356.000000 486.150000 ;
        RECT 351.000000 489.850000 356.000000 490.150000 ;
        RECT 401.000000 417.850000 406.000000 418.150000 ;
        RECT 401.000000 421.850000 406.000000 422.150000 ;
        RECT 401.000000 425.850000 406.000000 426.150000 ;
        RECT 401.000000 433.850000 406.000000 434.150000 ;
        RECT 401.000000 429.850000 406.000000 430.150000 ;
        RECT 401.000000 437.850000 406.000000 438.150000 ;
        RECT 401.000000 441.850000 406.000000 442.150000 ;
        RECT 401.000000 445.850000 406.000000 446.150000 ;
        RECT 401.000000 449.850000 406.000000 450.150000 ;
        RECT 401.000000 453.850000 406.000000 454.150000 ;
        RECT 401.000000 461.850000 406.000000 462.150000 ;
        RECT 401.000000 457.850000 406.000000 458.150000 ;
        RECT 401.000000 465.850000 406.000000 466.150000 ;
        RECT 401.000000 469.850000 406.000000 470.150000 ;
        RECT 401.000000 481.850000 406.000000 482.150000 ;
        RECT 401.000000 473.850000 406.000000 474.150000 ;
        RECT 401.000000 477.850000 406.000000 478.150000 ;
        RECT 401.000000 485.850000 406.000000 486.150000 ;
        RECT 401.000000 489.850000 406.000000 490.150000 ;
        RECT 451.000000 345.850000 456.000000 346.150000 ;
        RECT 451.000000 369.850000 456.000000 370.150000 ;
        RECT 451.000000 377.850000 456.000000 378.150000 ;
        RECT 451.000000 373.850000 456.000000 374.150000 ;
        RECT 501.000000 345.850000 506.000000 346.150000 ;
        RECT 501.000000 349.850000 506.000000 350.150000 ;
        RECT 501.000000 353.850000 506.000000 354.150000 ;
        RECT 501.000000 357.850000 506.000000 358.150000 ;
        RECT 501.000000 361.850000 506.000000 362.150000 ;
        RECT 501.000000 365.850000 506.000000 366.150000 ;
        RECT 501.000000 369.850000 506.000000 370.150000 ;
        RECT 501.000000 377.850000 506.000000 378.150000 ;
        RECT 501.000000 373.850000 506.000000 374.150000 ;
        RECT 451.000000 381.850000 456.000000 382.150000 ;
        RECT 451.000000 385.850000 456.000000 386.150000 ;
        RECT 451.000000 397.850000 456.000000 398.150000 ;
        RECT 451.000000 393.850000 456.000000 394.150000 ;
        RECT 451.000000 389.850000 456.000000 390.150000 ;
        RECT 501.000000 381.850000 506.000000 382.150000 ;
        RECT 501.000000 385.850000 506.000000 386.150000 ;
        RECT 501.000000 393.850000 506.000000 394.150000 ;
        RECT 501.000000 389.850000 506.000000 390.150000 ;
        RECT 501.000000 397.850000 506.000000 398.150000 ;
        RECT 501.000000 401.850000 506.000000 402.150000 ;
        RECT 501.000000 405.850000 506.000000 406.150000 ;
        RECT 501.000000 409.850000 506.000000 410.150000 ;
        RECT 501.000000 413.850000 506.000000 414.150000 ;
        RECT 551.000000 357.850000 556.000000 358.150000 ;
        RECT 551.000000 353.850000 556.000000 354.150000 ;
        RECT 551.000000 349.850000 556.000000 350.150000 ;
        RECT 551.000000 345.850000 556.000000 346.150000 ;
        RECT 551.000000 361.850000 556.000000 362.150000 ;
        RECT 551.000000 365.850000 556.000000 366.150000 ;
        RECT 551.000000 369.850000 556.000000 370.150000 ;
        RECT 551.000000 373.850000 556.000000 374.150000 ;
        RECT 551.000000 377.850000 556.000000 378.150000 ;
        RECT 551.000000 385.850000 556.000000 386.150000 ;
        RECT 551.000000 381.850000 556.000000 382.150000 ;
        RECT 551.000000 397.850000 556.000000 398.150000 ;
        RECT 551.000000 393.850000 556.000000 394.150000 ;
        RECT 551.000000 389.850000 556.000000 390.150000 ;
        RECT 551.000000 413.850000 556.000000 414.150000 ;
        RECT 551.000000 409.850000 556.000000 410.150000 ;
        RECT 551.000000 405.850000 556.000000 406.150000 ;
        RECT 551.000000 401.850000 556.000000 402.150000 ;
        RECT 451.000000 425.850000 456.000000 426.150000 ;
        RECT 451.000000 421.850000 456.000000 422.150000 ;
        RECT 451.000000 429.850000 456.000000 430.150000 ;
        RECT 451.000000 433.850000 456.000000 434.150000 ;
        RECT 451.000000 441.850000 456.000000 442.150000 ;
        RECT 451.000000 437.850000 456.000000 438.150000 ;
        RECT 451.000000 453.850000 456.000000 454.150000 ;
        RECT 451.000000 449.850000 456.000000 450.150000 ;
        RECT 451.000000 445.850000 456.000000 446.150000 ;
        RECT 501.000000 425.850000 506.000000 426.150000 ;
        RECT 501.000000 421.850000 506.000000 422.150000 ;
        RECT 501.000000 417.850000 506.000000 418.150000 ;
        RECT 501.000000 433.850000 506.000000 434.150000 ;
        RECT 501.000000 429.850000 506.000000 430.150000 ;
        RECT 501.000000 437.850000 506.000000 438.150000 ;
        RECT 501.000000 441.850000 506.000000 442.150000 ;
        RECT 501.000000 445.850000 506.000000 446.150000 ;
        RECT 501.000000 453.850000 506.000000 454.150000 ;
        RECT 501.000000 449.850000 506.000000 450.150000 ;
        RECT 451.000000 461.850000 456.000000 462.150000 ;
        RECT 451.000000 457.850000 456.000000 458.150000 ;
        RECT 451.000000 465.850000 456.000000 466.150000 ;
        RECT 451.000000 469.850000 456.000000 470.150000 ;
        RECT 451.000000 481.850000 456.000000 482.150000 ;
        RECT 451.000000 477.850000 456.000000 478.150000 ;
        RECT 451.000000 473.850000 456.000000 474.150000 ;
        RECT 451.000000 489.850000 456.000000 490.150000 ;
        RECT 451.000000 485.850000 456.000000 486.150000 ;
        RECT 501.000000 457.850000 506.000000 458.150000 ;
        RECT 501.000000 461.850000 506.000000 462.150000 ;
        RECT 501.000000 469.850000 506.000000 470.150000 ;
        RECT 501.000000 465.850000 506.000000 466.150000 ;
        RECT 501.000000 481.850000 506.000000 482.150000 ;
        RECT 501.000000 473.850000 506.000000 474.150000 ;
        RECT 501.000000 477.850000 506.000000 478.150000 ;
        RECT 501.000000 485.850000 506.000000 486.150000 ;
        RECT 501.000000 489.850000 506.000000 490.150000 ;
        RECT 551.000000 421.850000 556.000000 422.150000 ;
        RECT 551.000000 417.850000 556.000000 418.150000 ;
        RECT 551.000000 425.850000 556.000000 426.150000 ;
        RECT 551.000000 433.850000 556.000000 434.150000 ;
        RECT 551.000000 429.850000 556.000000 430.150000 ;
        RECT 551.000000 437.850000 556.000000 438.150000 ;
        RECT 551.000000 441.850000 556.000000 442.150000 ;
        RECT 551.000000 445.850000 556.000000 446.150000 ;
        RECT 551.000000 449.850000 556.000000 450.150000 ;
        RECT 551.000000 453.850000 556.000000 454.150000 ;
        RECT 551.000000 457.850000 556.000000 458.150000 ;
        RECT 551.000000 461.850000 556.000000 462.150000 ;
        RECT 551.000000 465.850000 556.000000 466.150000 ;
        RECT 551.000000 469.850000 556.000000 470.150000 ;
        RECT 551.000000 481.850000 556.000000 482.150000 ;
        RECT 551.000000 473.850000 556.000000 474.150000 ;
        RECT 551.000000 477.850000 556.000000 478.150000 ;
        RECT 551.000000 485.850000 556.000000 486.150000 ;
        RECT 551.000000 489.850000 556.000000 490.150000 ;
        RECT 301.000000 497.850000 306.000000 498.150000 ;
        RECT 301.000000 493.850000 306.000000 494.150000 ;
        RECT 301.000000 501.850000 306.000000 502.150000 ;
        RECT 301.000000 505.850000 306.000000 506.150000 ;
        RECT 301.000000 517.850000 306.000000 518.150000 ;
        RECT 301.000000 513.850000 306.000000 514.150000 ;
        RECT 301.000000 509.850000 306.000000 510.150000 ;
        RECT 351.000000 497.850000 356.000000 498.150000 ;
        RECT 351.000000 493.850000 356.000000 494.150000 ;
        RECT 351.000000 501.850000 356.000000 502.150000 ;
        RECT 351.000000 505.850000 356.000000 506.150000 ;
        RECT 351.000000 509.850000 356.000000 510.150000 ;
        RECT 351.000000 513.850000 356.000000 514.150000 ;
        RECT 351.000000 517.850000 356.000000 518.150000 ;
        RECT 351.000000 521.850000 356.000000 522.150000 ;
        RECT 351.000000 525.850000 356.000000 526.150000 ;
        RECT 351.000000 529.850000 356.000000 530.150000 ;
        RECT 351.000000 533.850000 356.000000 534.150000 ;
        RECT 351.000000 545.850000 356.000000 546.150000 ;
        RECT 351.000000 541.850000 356.000000 542.150000 ;
        RECT 351.000000 537.850000 356.000000 538.150000 ;
        RECT 351.000000 561.850000 356.000000 562.150000 ;
        RECT 351.000000 557.850000 356.000000 558.150000 ;
        RECT 351.000000 553.850000 356.000000 554.150000 ;
        RECT 351.000000 549.850000 356.000000 550.150000 ;
        RECT 385.000000 505.850000 395.000000 506.150000 ;
        RECT 385.000000 501.850000 395.000000 502.150000 ;
        RECT 385.000000 493.850000 395.000000 494.150000 ;
        RECT 385.000000 497.850000 395.000000 498.150000 ;
        RECT 401.000000 497.850000 406.000000 498.150000 ;
        RECT 401.000000 493.850000 406.000000 494.150000 ;
        RECT 401.000000 501.850000 406.000000 502.150000 ;
        RECT 385.000000 509.850000 395.000000 510.150000 ;
        RECT 385.000000 513.850000 395.000000 514.150000 ;
        RECT 385.000000 517.850000 395.000000 518.150000 ;
        RECT 385.000000 521.850000 395.000000 522.150000 ;
        RECT 385.000000 525.850000 395.000000 526.150000 ;
        RECT 385.000000 545.850000 395.000000 546.150000 ;
        RECT 385.000000 541.850000 395.000000 542.150000 ;
        RECT 385.000000 537.850000 395.000000 538.150000 ;
        RECT 385.000000 533.850000 395.000000 534.150000 ;
        RECT 385.000000 529.850000 395.000000 530.150000 ;
        RECT 385.000000 561.850000 395.000000 562.150000 ;
        RECT 385.000000 557.850000 395.000000 558.150000 ;
        RECT 385.000000 553.850000 395.000000 554.150000 ;
        RECT 385.000000 549.850000 395.000000 550.150000 ;
        RECT 351.000000 565.850000 356.000000 566.150000 ;
        RECT 351.000000 569.850000 356.000000 570.150000 ;
        RECT 351.000000 573.850000 356.000000 574.150000 ;
        RECT 351.000000 577.850000 356.000000 578.150000 ;
        RECT 351.000000 581.850000 356.000000 582.150000 ;
        RECT 351.000000 601.850000 356.000000 602.150000 ;
        RECT 351.000000 597.850000 356.000000 598.150000 ;
        RECT 351.000000 593.850000 356.000000 594.150000 ;
        RECT 351.000000 589.850000 356.000000 590.150000 ;
        RECT 351.000000 585.850000 356.000000 586.150000 ;
        RECT 351.000000 609.850000 356.000000 610.150000 ;
        RECT 351.000000 605.850000 356.000000 606.150000 ;
        RECT 351.000000 613.850000 356.000000 614.150000 ;
        RECT 351.000000 617.850000 356.000000 618.150000 ;
        RECT 351.000000 621.850000 356.000000 622.150000 ;
        RECT 351.000000 625.850000 356.000000 626.150000 ;
        RECT 351.000000 629.850000 356.000000 630.150000 ;
        RECT 351.000000 633.850000 356.000000 634.150000 ;
        RECT 351.000000 637.850000 356.000000 638.150000 ;
        RECT 385.000000 581.850000 395.000000 582.150000 ;
        RECT 385.000000 565.850000 395.000000 566.150000 ;
        RECT 385.000000 569.850000 395.000000 570.150000 ;
        RECT 385.000000 573.850000 395.000000 574.150000 ;
        RECT 385.000000 577.850000 395.000000 578.150000 ;
        RECT 385.000000 601.850000 395.000000 602.150000 ;
        RECT 385.000000 597.850000 395.000000 598.150000 ;
        RECT 385.000000 593.850000 395.000000 594.150000 ;
        RECT 385.000000 589.850000 395.000000 590.150000 ;
        RECT 385.000000 585.850000 395.000000 586.150000 ;
        RECT 385.000000 617.850000 395.000000 618.150000 ;
        RECT 385.000000 613.850000 395.000000 614.150000 ;
        RECT 385.000000 609.850000 395.000000 610.150000 ;
        RECT 385.000000 605.850000 395.000000 606.150000 ;
        RECT 385.000000 637.850000 395.000000 638.150000 ;
        RECT 385.000000 633.850000 395.000000 634.150000 ;
        RECT 385.000000 629.850000 395.000000 630.150000 ;
        RECT 385.000000 625.850000 395.000000 626.150000 ;
        RECT 385.000000 621.850000 395.000000 622.150000 ;
        RECT 451.000000 493.850000 456.000000 494.150000 ;
        RECT 451.000000 497.850000 456.000000 498.150000 ;
        RECT 451.000000 501.850000 456.000000 502.150000 ;
        RECT 501.000000 493.850000 506.000000 494.150000 ;
        RECT 501.000000 497.850000 506.000000 498.150000 ;
        RECT 501.000000 501.850000 506.000000 502.150000 ;
        RECT 551.000000 493.850000 556.000000 494.150000 ;
        RECT 551.000000 497.850000 556.000000 498.150000 ;
        RECT 551.000000 501.850000 556.000000 502.150000 ;
        RECT 351.000000 657.850000 356.000000 658.150000 ;
        RECT 351.000000 641.850000 356.000000 642.150000 ;
        RECT 351.000000 645.850000 356.000000 646.150000 ;
        RECT 351.000000 649.850000 356.000000 650.150000 ;
        RECT 351.000000 653.850000 356.000000 654.150000 ;
        RECT 351.000000 673.850000 356.000000 674.150000 ;
        RECT 351.000000 669.850000 356.000000 670.150000 ;
        RECT 351.000000 665.850000 356.000000 666.150000 ;
        RECT 351.000000 661.850000 356.000000 662.150000 ;
        RECT 301.000000 681.850000 306.000000 682.150000 ;
        RECT 301.000000 677.850000 306.000000 678.150000 ;
        RECT 351.000000 677.850000 356.000000 678.150000 ;
        RECT 351.000000 681.850000 356.000000 682.150000 ;
        RECT 385.000000 657.850000 395.000000 658.150000 ;
        RECT 401.000000 657.850000 406.000000 658.150000 ;
        RECT 385.000000 641.850000 395.000000 642.150000 ;
        RECT 385.000000 645.850000 395.000000 646.150000 ;
        RECT 385.000000 649.850000 395.000000 650.150000 ;
        RECT 385.000000 653.850000 395.000000 654.150000 ;
        RECT 385.000000 673.850000 395.000000 674.150000 ;
        RECT 385.000000 669.850000 395.000000 670.150000 ;
        RECT 385.000000 665.850000 395.000000 666.150000 ;
        RECT 385.000000 661.850000 395.000000 662.150000 ;
        RECT 401.000000 661.850000 406.000000 662.150000 ;
        RECT 401.000000 665.850000 406.000000 666.150000 ;
        RECT 401.000000 669.850000 406.000000 670.150000 ;
        RECT 401.000000 673.850000 406.000000 674.150000 ;
        RECT 401.000000 677.850000 406.000000 678.150000 ;
        RECT 385.000000 677.850000 395.000000 678.150000 ;
        RECT 401.000000 681.850000 406.000000 682.150000 ;
        RECT 385.000000 681.850000 395.000000 682.150000 ;
        RECT 451.000000 657.850000 456.000000 658.150000 ;
        RECT 451.000000 661.850000 456.000000 662.150000 ;
        RECT 451.000000 665.850000 456.000000 666.150000 ;
        RECT 451.000000 669.850000 456.000000 670.150000 ;
        RECT 451.000000 673.850000 456.000000 674.150000 ;
        RECT 501.000000 657.850000 506.000000 658.150000 ;
        RECT 501.000000 661.850000 506.000000 662.150000 ;
        RECT 501.000000 665.850000 506.000000 666.150000 ;
        RECT 501.000000 673.850000 506.000000 674.150000 ;
        RECT 501.000000 669.850000 506.000000 670.150000 ;
        RECT 451.000000 677.850000 456.000000 678.150000 ;
        RECT 451.000000 681.850000 456.000000 682.150000 ;
        RECT 501.000000 677.850000 506.000000 678.150000 ;
        RECT 501.000000 681.850000 506.000000 682.150000 ;
        RECT 551.000000 673.850000 556.000000 674.150000 ;
        RECT 551.000000 657.850000 556.000000 658.150000 ;
        RECT 551.000000 661.850000 556.000000 662.150000 ;
        RECT 551.000000 665.850000 556.000000 666.150000 ;
        RECT 551.000000 669.850000 556.000000 670.150000 ;
        RECT 551.000000 681.850000 556.000000 682.150000 ;
        RECT 551.000000 677.850000 556.000000 678.150000 ;
        RECT 735.000000 433.850000 745.000000 434.150000 ;
        RECT 735.000000 441.850000 745.000000 442.150000 ;
        RECT 735.000000 437.850000 745.000000 438.150000 ;
        RECT 735.000000 445.850000 745.000000 446.150000 ;
        RECT 735.000000 449.850000 745.000000 450.150000 ;
        RECT 735.000000 453.850000 745.000000 454.150000 ;
        RECT 735.000000 457.850000 745.000000 458.150000 ;
        RECT 735.000000 461.850000 745.000000 462.150000 ;
        RECT 735.000000 465.850000 745.000000 466.150000 ;
        RECT 735.000000 469.850000 745.000000 470.150000 ;
        RECT 735.000000 481.850000 745.000000 482.150000 ;
        RECT 735.000000 473.850000 745.000000 474.150000 ;
        RECT 735.000000 477.850000 745.000000 478.150000 ;
        RECT 735.000000 485.850000 745.000000 486.150000 ;
        RECT 735.000000 489.850000 745.000000 490.150000 ;
        RECT 601.000000 357.850000 606.000000 358.150000 ;
        RECT 601.000000 353.850000 606.000000 354.150000 ;
        RECT 601.000000 345.850000 606.000000 346.150000 ;
        RECT 601.000000 349.850000 606.000000 350.150000 ;
        RECT 601.000000 361.850000 606.000000 362.150000 ;
        RECT 601.000000 365.850000 606.000000 366.150000 ;
        RECT 601.000000 369.850000 606.000000 370.150000 ;
        RECT 601.000000 373.850000 606.000000 374.150000 ;
        RECT 601.000000 377.850000 606.000000 378.150000 ;
        RECT 651.000000 349.850000 656.000000 350.150000 ;
        RECT 651.000000 345.850000 656.000000 346.150000 ;
        RECT 651.000000 353.850000 656.000000 354.150000 ;
        RECT 651.000000 357.850000 656.000000 358.150000 ;
        RECT 651.000000 361.850000 656.000000 362.150000 ;
        RECT 651.000000 365.850000 656.000000 366.150000 ;
        RECT 651.000000 369.850000 656.000000 370.150000 ;
        RECT 651.000000 373.850000 656.000000 374.150000 ;
        RECT 651.000000 377.850000 656.000000 378.150000 ;
        RECT 601.000000 385.850000 606.000000 386.150000 ;
        RECT 601.000000 381.850000 606.000000 382.150000 ;
        RECT 601.000000 397.850000 606.000000 398.150000 ;
        RECT 601.000000 389.850000 606.000000 390.150000 ;
        RECT 601.000000 393.850000 606.000000 394.150000 ;
        RECT 601.000000 405.850000 606.000000 406.150000 ;
        RECT 601.000000 401.850000 606.000000 402.150000 ;
        RECT 601.000000 413.850000 606.000000 414.150000 ;
        RECT 601.000000 409.850000 606.000000 410.150000 ;
        RECT 651.000000 381.850000 656.000000 382.150000 ;
        RECT 651.000000 385.850000 656.000000 386.150000 ;
        RECT 651.000000 393.850000 656.000000 394.150000 ;
        RECT 651.000000 389.850000 656.000000 390.150000 ;
        RECT 651.000000 397.850000 656.000000 398.150000 ;
        RECT 651.000000 401.850000 656.000000 402.150000 ;
        RECT 651.000000 405.850000 656.000000 406.150000 ;
        RECT 651.000000 409.850000 656.000000 410.150000 ;
        RECT 651.000000 413.850000 656.000000 414.150000 ;
        RECT 701.000000 357.850000 706.000000 358.150000 ;
        RECT 701.000000 353.850000 706.000000 354.150000 ;
        RECT 701.000000 349.850000 706.000000 350.150000 ;
        RECT 701.000000 345.850000 706.000000 346.150000 ;
        RECT 701.000000 361.850000 706.000000 362.150000 ;
        RECT 701.000000 365.850000 706.000000 366.150000 ;
        RECT 701.000000 369.850000 706.000000 370.150000 ;
        RECT 701.000000 373.850000 706.000000 374.150000 ;
        RECT 701.000000 377.850000 706.000000 378.150000 ;
        RECT 701.000000 385.850000 706.000000 386.150000 ;
        RECT 701.000000 381.850000 706.000000 382.150000 ;
        RECT 701.000000 397.850000 706.000000 398.150000 ;
        RECT 701.000000 393.850000 706.000000 394.150000 ;
        RECT 701.000000 389.850000 706.000000 390.150000 ;
        RECT 701.000000 413.850000 706.000000 414.150000 ;
        RECT 701.000000 409.850000 706.000000 410.150000 ;
        RECT 701.000000 405.850000 706.000000 406.150000 ;
        RECT 701.000000 401.850000 706.000000 402.150000 ;
        RECT 601.000000 417.850000 606.000000 418.150000 ;
        RECT 601.000000 421.850000 606.000000 422.150000 ;
        RECT 601.000000 425.850000 606.000000 426.150000 ;
        RECT 601.000000 429.850000 606.000000 430.150000 ;
        RECT 601.000000 433.850000 606.000000 434.150000 ;
        RECT 601.000000 441.850000 606.000000 442.150000 ;
        RECT 601.000000 437.850000 606.000000 438.150000 ;
        RECT 601.000000 453.850000 606.000000 454.150000 ;
        RECT 601.000000 449.850000 606.000000 450.150000 ;
        RECT 601.000000 445.850000 606.000000 446.150000 ;
        RECT 651.000000 417.850000 656.000000 418.150000 ;
        RECT 651.000000 425.850000 656.000000 426.150000 ;
        RECT 651.000000 421.850000 656.000000 422.150000 ;
        RECT 651.000000 429.850000 656.000000 430.150000 ;
        RECT 651.000000 433.850000 656.000000 434.150000 ;
        RECT 651.000000 437.850000 656.000000 438.150000 ;
        RECT 651.000000 441.850000 656.000000 442.150000 ;
        RECT 651.000000 445.850000 656.000000 446.150000 ;
        RECT 651.000000 449.850000 656.000000 450.150000 ;
        RECT 651.000000 453.850000 656.000000 454.150000 ;
        RECT 601.000000 461.850000 606.000000 462.150000 ;
        RECT 601.000000 457.850000 606.000000 458.150000 ;
        RECT 601.000000 465.850000 606.000000 466.150000 ;
        RECT 601.000000 469.850000 606.000000 470.150000 ;
        RECT 601.000000 481.850000 606.000000 482.150000 ;
        RECT 601.000000 477.850000 606.000000 478.150000 ;
        RECT 601.000000 473.850000 606.000000 474.150000 ;
        RECT 601.000000 489.850000 606.000000 490.150000 ;
        RECT 601.000000 485.850000 606.000000 486.150000 ;
        RECT 651.000000 457.850000 656.000000 458.150000 ;
        RECT 651.000000 461.850000 656.000000 462.150000 ;
        RECT 651.000000 469.850000 656.000000 470.150000 ;
        RECT 651.000000 465.850000 656.000000 466.150000 ;
        RECT 651.000000 481.850000 656.000000 482.150000 ;
        RECT 651.000000 477.850000 656.000000 478.150000 ;
        RECT 651.000000 473.850000 656.000000 474.150000 ;
        RECT 651.000000 489.850000 656.000000 490.150000 ;
        RECT 651.000000 485.850000 656.000000 486.150000 ;
        RECT 701.000000 417.850000 706.000000 418.150000 ;
        RECT 701.000000 421.850000 706.000000 422.150000 ;
        RECT 701.000000 425.850000 706.000000 426.150000 ;
        RECT 701.000000 433.850000 706.000000 434.150000 ;
        RECT 701.000000 429.850000 706.000000 430.150000 ;
        RECT 701.000000 437.850000 706.000000 438.150000 ;
        RECT 701.000000 441.850000 706.000000 442.150000 ;
        RECT 701.000000 445.850000 706.000000 446.150000 ;
        RECT 701.000000 449.850000 706.000000 450.150000 ;
        RECT 701.000000 453.850000 706.000000 454.150000 ;
        RECT 701.000000 457.850000 706.000000 458.150000 ;
        RECT 701.000000 461.850000 706.000000 462.150000 ;
        RECT 701.000000 465.850000 706.000000 466.150000 ;
        RECT 701.000000 469.850000 706.000000 470.150000 ;
        RECT 701.000000 481.850000 706.000000 482.150000 ;
        RECT 701.000000 473.850000 706.000000 474.150000 ;
        RECT 701.000000 477.850000 706.000000 478.150000 ;
        RECT 701.000000 485.850000 706.000000 486.150000 ;
        RECT 701.000000 489.850000 706.000000 490.150000 ;
        RECT 751.000000 357.850000 756.000000 358.150000 ;
        RECT 751.000000 353.850000 756.000000 354.150000 ;
        RECT 751.000000 349.850000 756.000000 350.150000 ;
        RECT 751.000000 345.850000 756.000000 346.150000 ;
        RECT 751.000000 361.850000 756.000000 362.150000 ;
        RECT 751.000000 365.850000 756.000000 366.150000 ;
        RECT 751.000000 369.850000 756.000000 370.150000 ;
        RECT 751.000000 373.850000 756.000000 374.150000 ;
        RECT 751.000000 377.850000 756.000000 378.150000 ;
        RECT 801.000000 345.850000 806.000000 346.150000 ;
        RECT 801.000000 349.850000 806.000000 350.150000 ;
        RECT 801.000000 353.850000 806.000000 354.150000 ;
        RECT 801.000000 357.850000 806.000000 358.150000 ;
        RECT 801.000000 361.850000 806.000000 362.150000 ;
        RECT 801.000000 365.850000 806.000000 366.150000 ;
        RECT 801.000000 369.850000 806.000000 370.150000 ;
        RECT 801.000000 377.850000 806.000000 378.150000 ;
        RECT 801.000000 373.850000 806.000000 374.150000 ;
        RECT 751.000000 385.850000 756.000000 386.150000 ;
        RECT 751.000000 381.850000 756.000000 382.150000 ;
        RECT 751.000000 393.850000 756.000000 394.150000 ;
        RECT 751.000000 389.850000 756.000000 390.150000 ;
        RECT 751.000000 397.850000 756.000000 398.150000 ;
        RECT 751.000000 401.850000 756.000000 402.150000 ;
        RECT 751.000000 405.850000 756.000000 406.150000 ;
        RECT 751.000000 413.850000 756.000000 414.150000 ;
        RECT 751.000000 409.850000 756.000000 410.150000 ;
        RECT 801.000000 385.850000 806.000000 386.150000 ;
        RECT 801.000000 381.850000 806.000000 382.150000 ;
        RECT 801.000000 393.850000 806.000000 394.150000 ;
        RECT 801.000000 389.850000 806.000000 390.150000 ;
        RECT 801.000000 397.850000 806.000000 398.150000 ;
        RECT 801.000000 401.850000 806.000000 402.150000 ;
        RECT 801.000000 405.850000 806.000000 406.150000 ;
        RECT 801.000000 413.850000 806.000000 414.150000 ;
        RECT 801.000000 409.850000 806.000000 410.150000 ;
        RECT 851.000000 357.850000 856.000000 358.150000 ;
        RECT 851.000000 353.850000 856.000000 354.150000 ;
        RECT 851.000000 349.850000 856.000000 350.150000 ;
        RECT 851.000000 345.850000 856.000000 346.150000 ;
        RECT 851.000000 361.850000 856.000000 362.150000 ;
        RECT 851.000000 365.850000 856.000000 366.150000 ;
        RECT 851.000000 369.850000 856.000000 370.150000 ;
        RECT 851.000000 373.850000 856.000000 374.150000 ;
        RECT 851.000000 377.850000 856.000000 378.150000 ;
        RECT 851.000000 385.850000 856.000000 386.150000 ;
        RECT 851.000000 381.850000 856.000000 382.150000 ;
        RECT 851.000000 397.850000 856.000000 398.150000 ;
        RECT 851.000000 393.850000 856.000000 394.150000 ;
        RECT 851.000000 389.850000 856.000000 390.150000 ;
        RECT 851.000000 413.850000 856.000000 414.150000 ;
        RECT 851.000000 409.850000 856.000000 410.150000 ;
        RECT 851.000000 405.850000 856.000000 406.150000 ;
        RECT 851.000000 401.850000 856.000000 402.150000 ;
        RECT 751.000000 417.850000 756.000000 418.150000 ;
        RECT 751.000000 421.850000 756.000000 422.150000 ;
        RECT 751.000000 425.850000 756.000000 426.150000 ;
        RECT 751.000000 429.850000 756.000000 430.150000 ;
        RECT 751.000000 433.850000 756.000000 434.150000 ;
        RECT 751.000000 437.850000 756.000000 438.150000 ;
        RECT 751.000000 441.850000 756.000000 442.150000 ;
        RECT 801.000000 417.850000 806.000000 418.150000 ;
        RECT 801.000000 421.850000 806.000000 422.150000 ;
        RECT 801.000000 425.850000 806.000000 426.150000 ;
        RECT 801.000000 429.850000 806.000000 430.150000 ;
        RECT 801.000000 433.850000 806.000000 434.150000 ;
        RECT 801.000000 437.850000 806.000000 438.150000 ;
        RECT 801.000000 441.850000 806.000000 442.150000 ;
        RECT 851.000000 429.850000 856.000000 430.150000 ;
        RECT 851.000000 425.850000 856.000000 426.150000 ;
        RECT 851.000000 421.850000 856.000000 422.150000 ;
        RECT 851.000000 417.850000 856.000000 418.150000 ;
        RECT 851.000000 433.850000 856.000000 434.150000 ;
        RECT 851.000000 441.850000 856.000000 442.150000 ;
        RECT 851.000000 437.850000 856.000000 438.150000 ;
        RECT 735.000000 501.850000 745.000000 502.150000 ;
        RECT 735.000000 497.850000 745.000000 498.150000 ;
        RECT 735.000000 493.850000 745.000000 494.150000 ;
        RECT 601.000000 501.850000 606.000000 502.150000 ;
        RECT 601.000000 497.850000 606.000000 498.150000 ;
        RECT 601.000000 493.850000 606.000000 494.150000 ;
        RECT 651.000000 497.850000 656.000000 498.150000 ;
        RECT 651.000000 493.850000 656.000000 494.150000 ;
        RECT 651.000000 501.850000 656.000000 502.150000 ;
        RECT 701.000000 493.850000 706.000000 494.150000 ;
        RECT 701.000000 497.850000 706.000000 498.150000 ;
        RECT 701.000000 501.850000 706.000000 502.150000 ;
        RECT 901.000000 357.850000 906.000000 358.150000 ;
        RECT 901.000000 353.850000 906.000000 354.150000 ;
        RECT 901.000000 349.850000 906.000000 350.150000 ;
        RECT 901.000000 345.850000 906.000000 346.150000 ;
        RECT 901.000000 361.850000 906.000000 362.150000 ;
        RECT 901.000000 365.850000 906.000000 366.150000 ;
        RECT 901.000000 369.850000 906.000000 370.150000 ;
        RECT 901.000000 373.850000 906.000000 374.150000 ;
        RECT 901.000000 377.850000 906.000000 378.150000 ;
        RECT 951.000000 345.850000 956.000000 346.150000 ;
        RECT 951.000000 349.850000 956.000000 350.150000 ;
        RECT 951.000000 353.850000 956.000000 354.150000 ;
        RECT 951.000000 357.850000 956.000000 358.150000 ;
        RECT 951.000000 361.850000 956.000000 362.150000 ;
        RECT 951.000000 365.850000 956.000000 366.150000 ;
        RECT 951.000000 369.850000 956.000000 370.150000 ;
        RECT 951.000000 373.850000 956.000000 374.150000 ;
        RECT 951.000000 377.850000 956.000000 378.150000 ;
        RECT 901.000000 385.850000 906.000000 386.150000 ;
        RECT 901.000000 381.850000 906.000000 382.150000 ;
        RECT 901.000000 393.850000 906.000000 394.150000 ;
        RECT 901.000000 389.850000 906.000000 390.150000 ;
        RECT 901.000000 397.850000 906.000000 398.150000 ;
        RECT 901.000000 401.850000 906.000000 402.150000 ;
        RECT 901.000000 405.850000 906.000000 406.150000 ;
        RECT 901.000000 413.850000 906.000000 414.150000 ;
        RECT 901.000000 409.850000 906.000000 410.150000 ;
        RECT 951.000000 385.850000 956.000000 386.150000 ;
        RECT 951.000000 381.850000 956.000000 382.150000 ;
        RECT 951.000000 389.850000 956.000000 390.150000 ;
        RECT 951.000000 393.850000 956.000000 394.150000 ;
        RECT 951.000000 397.850000 956.000000 398.150000 ;
        RECT 951.000000 405.850000 956.000000 406.150000 ;
        RECT 951.000000 401.850000 956.000000 402.150000 ;
        RECT 951.000000 413.850000 956.000000 414.150000 ;
        RECT 951.000000 409.850000 956.000000 410.150000 ;
        RECT 1001.000000 349.850000 1006.000000 350.150000 ;
        RECT 1001.000000 345.850000 1006.000000 346.150000 ;
        RECT 1001.000000 353.850000 1006.000000 354.150000 ;
        RECT 1001.000000 357.850000 1006.000000 358.150000 ;
        RECT 1001.000000 361.850000 1006.000000 362.150000 ;
        RECT 1001.000000 365.850000 1006.000000 366.150000 ;
        RECT 1001.000000 369.850000 1006.000000 370.150000 ;
        RECT 1001.000000 377.850000 1006.000000 378.150000 ;
        RECT 1001.000000 373.850000 1006.000000 374.150000 ;
        RECT 1001.000000 385.850000 1006.000000 386.150000 ;
        RECT 1001.000000 381.850000 1006.000000 382.150000 ;
        RECT 1001.000000 393.850000 1006.000000 394.150000 ;
        RECT 1001.000000 389.850000 1006.000000 390.150000 ;
        RECT 1001.000000 397.850000 1006.000000 398.150000 ;
        RECT 1001.000000 405.850000 1006.000000 406.150000 ;
        RECT 1001.000000 401.850000 1006.000000 402.150000 ;
        RECT 1001.000000 413.850000 1006.000000 414.150000 ;
        RECT 1001.000000 409.850000 1006.000000 410.150000 ;
        RECT 901.000000 417.850000 906.000000 418.150000 ;
        RECT 901.000000 421.850000 906.000000 422.150000 ;
        RECT 901.000000 425.850000 906.000000 426.150000 ;
        RECT 901.000000 429.850000 906.000000 430.150000 ;
        RECT 901.000000 433.850000 906.000000 434.150000 ;
        RECT 901.000000 437.850000 906.000000 438.150000 ;
        RECT 901.000000 441.850000 906.000000 442.150000 ;
        RECT 951.000000 417.850000 956.000000 418.150000 ;
        RECT 951.000000 421.850000 956.000000 422.150000 ;
        RECT 951.000000 425.850000 956.000000 426.150000 ;
        RECT 951.000000 429.850000 956.000000 430.150000 ;
        RECT 951.000000 433.850000 956.000000 434.150000 ;
        RECT 951.000000 441.850000 956.000000 442.150000 ;
        RECT 951.000000 437.850000 956.000000 438.150000 ;
        RECT 1001.000000 425.850000 1006.000000 426.150000 ;
        RECT 1001.000000 421.850000 1006.000000 422.150000 ;
        RECT 1001.000000 417.850000 1006.000000 418.150000 ;
        RECT 1001.000000 429.850000 1006.000000 430.150000 ;
        RECT 1001.000000 433.850000 1006.000000 434.150000 ;
        RECT 1001.000000 437.850000 1006.000000 438.150000 ;
        RECT 1001.000000 441.850000 1006.000000 442.150000 ;
        RECT 1051.000000 357.850000 1056.000000 358.150000 ;
        RECT 1051.000000 353.850000 1056.000000 354.150000 ;
        RECT 1051.000000 349.850000 1056.000000 350.150000 ;
        RECT 1051.000000 345.850000 1056.000000 346.150000 ;
        RECT 1051.000000 361.850000 1056.000000 362.150000 ;
        RECT 1051.000000 365.850000 1056.000000 366.150000 ;
        RECT 1051.000000 369.850000 1056.000000 370.150000 ;
        RECT 1051.000000 373.850000 1056.000000 374.150000 ;
        RECT 1051.000000 377.850000 1056.000000 378.150000 ;
        RECT 1101.000000 345.850000 1106.000000 346.150000 ;
        RECT 1101.000000 349.850000 1106.000000 350.150000 ;
        RECT 1101.000000 353.850000 1106.000000 354.150000 ;
        RECT 1101.000000 357.850000 1106.000000 358.150000 ;
        RECT 1101.000000 361.850000 1106.000000 362.150000 ;
        RECT 1101.000000 365.850000 1106.000000 366.150000 ;
        RECT 1101.000000 369.850000 1106.000000 370.150000 ;
        RECT 1101.000000 373.850000 1106.000000 374.150000 ;
        RECT 1101.000000 377.850000 1106.000000 378.150000 ;
        RECT 1051.000000 385.850000 1056.000000 386.150000 ;
        RECT 1051.000000 381.850000 1056.000000 382.150000 ;
        RECT 1051.000000 393.850000 1056.000000 394.150000 ;
        RECT 1051.000000 389.850000 1056.000000 390.150000 ;
        RECT 1051.000000 397.850000 1056.000000 398.150000 ;
        RECT 1051.000000 401.850000 1056.000000 402.150000 ;
        RECT 1051.000000 405.850000 1056.000000 406.150000 ;
        RECT 1051.000000 413.850000 1056.000000 414.150000 ;
        RECT 1051.000000 409.850000 1056.000000 410.150000 ;
        RECT 1101.000000 385.850000 1106.000000 386.150000 ;
        RECT 1101.000000 381.850000 1106.000000 382.150000 ;
        RECT 1101.000000 389.850000 1106.000000 390.150000 ;
        RECT 1101.000000 393.850000 1106.000000 394.150000 ;
        RECT 1101.000000 397.850000 1106.000000 398.150000 ;
        RECT 1101.000000 405.850000 1106.000000 406.150000 ;
        RECT 1101.000000 401.850000 1106.000000 402.150000 ;
        RECT 1101.000000 413.850000 1106.000000 414.150000 ;
        RECT 1101.000000 409.850000 1106.000000 410.150000 ;
        RECT 1151.000000 357.850000 1156.000000 358.150000 ;
        RECT 1151.000000 353.850000 1156.000000 354.150000 ;
        RECT 1151.000000 349.850000 1156.000000 350.150000 ;
        RECT 1151.000000 345.850000 1156.000000 346.150000 ;
        RECT 1172.000000 357.850000 1182.000000 358.150000 ;
        RECT 1172.000000 349.850000 1182.000000 350.150000 ;
        RECT 1172.000000 345.850000 1182.000000 346.150000 ;
        RECT 1172.000000 353.850000 1182.000000 354.150000 ;
        RECT 1151.000000 365.850000 1156.000000 366.150000 ;
        RECT 1151.000000 361.850000 1156.000000 362.150000 ;
        RECT 1151.000000 369.850000 1156.000000 370.150000 ;
        RECT 1151.000000 373.850000 1156.000000 374.150000 ;
        RECT 1151.000000 377.850000 1156.000000 378.150000 ;
        RECT 1172.000000 369.850000 1182.000000 370.150000 ;
        RECT 1172.000000 365.850000 1182.000000 366.150000 ;
        RECT 1172.000000 361.850000 1182.000000 362.150000 ;
        RECT 1172.000000 373.850000 1182.000000 374.150000 ;
        RECT 1172.000000 377.850000 1182.000000 378.150000 ;
        RECT 1151.000000 385.850000 1156.000000 386.150000 ;
        RECT 1151.000000 381.850000 1156.000000 382.150000 ;
        RECT 1151.000000 389.850000 1156.000000 390.150000 ;
        RECT 1151.000000 393.850000 1156.000000 394.150000 ;
        RECT 1151.000000 397.850000 1156.000000 398.150000 ;
        RECT 1172.000000 385.850000 1182.000000 386.150000 ;
        RECT 1172.000000 381.850000 1182.000000 382.150000 ;
        RECT 1172.000000 389.850000 1182.000000 390.150000 ;
        RECT 1172.000000 393.850000 1182.000000 394.150000 ;
        RECT 1172.000000 397.850000 1182.000000 398.150000 ;
        RECT 1151.000000 405.850000 1156.000000 406.150000 ;
        RECT 1151.000000 401.850000 1156.000000 402.150000 ;
        RECT 1151.000000 409.850000 1156.000000 410.150000 ;
        RECT 1151.000000 413.850000 1156.000000 414.150000 ;
        RECT 1172.000000 405.850000 1182.000000 406.150000 ;
        RECT 1172.000000 401.850000 1182.000000 402.150000 ;
        RECT 1172.000000 409.850000 1182.000000 410.150000 ;
        RECT 1172.000000 413.850000 1182.000000 414.150000 ;
        RECT 1051.000000 417.850000 1056.000000 418.150000 ;
        RECT 1051.000000 421.850000 1056.000000 422.150000 ;
        RECT 1051.000000 425.850000 1056.000000 426.150000 ;
        RECT 1051.000000 429.850000 1056.000000 430.150000 ;
        RECT 1051.000000 433.850000 1056.000000 434.150000 ;
        RECT 1051.000000 437.850000 1056.000000 438.150000 ;
        RECT 1051.000000 441.850000 1056.000000 442.150000 ;
        RECT 1101.000000 433.850000 1106.000000 434.150000 ;
        RECT 1101.000000 429.850000 1106.000000 430.150000 ;
        RECT 1101.000000 425.850000 1106.000000 426.150000 ;
        RECT 1101.000000 421.850000 1106.000000 422.150000 ;
        RECT 1101.000000 417.850000 1106.000000 418.150000 ;
        RECT 1101.000000 441.850000 1106.000000 442.150000 ;
        RECT 1101.000000 437.850000 1106.000000 438.150000 ;
        RECT 1151.000000 417.850000 1156.000000 418.150000 ;
        RECT 1151.000000 421.850000 1156.000000 422.150000 ;
        RECT 1151.000000 425.850000 1156.000000 426.150000 ;
        RECT 1151.000000 429.850000 1156.000000 430.150000 ;
        RECT 1151.000000 433.850000 1156.000000 434.150000 ;
        RECT 1172.000000 417.850000 1182.000000 418.150000 ;
        RECT 1172.000000 421.850000 1182.000000 422.150000 ;
        RECT 1172.000000 425.850000 1182.000000 426.150000 ;
        RECT 1172.000000 429.850000 1182.000000 430.150000 ;
        RECT 1172.000000 433.850000 1182.000000 434.150000 ;
        RECT 1151.000000 437.850000 1156.000000 438.150000 ;
        RECT 1151.000000 441.850000 1156.000000 442.150000 ;
        RECT 1151.000000 453.850000 1156.000000 454.150000 ;
        RECT 1151.000000 449.850000 1156.000000 450.150000 ;
        RECT 1151.000000 445.850000 1156.000000 446.150000 ;
        RECT 1172.000000 437.850000 1182.000000 438.150000 ;
        RECT 1172.000000 441.850000 1182.000000 442.150000 ;
        RECT 1151.000000 461.850000 1156.000000 462.150000 ;
        RECT 1151.000000 457.850000 1156.000000 458.150000 ;
        RECT 1151.000000 465.850000 1156.000000 466.150000 ;
        RECT 1151.000000 469.850000 1156.000000 470.150000 ;
        RECT 1151.000000 481.850000 1156.000000 482.150000 ;
        RECT 1151.000000 477.850000 1156.000000 478.150000 ;
        RECT 1151.000000 473.850000 1156.000000 474.150000 ;
        RECT 1151.000000 489.850000 1156.000000 490.150000 ;
        RECT 1151.000000 485.850000 1156.000000 486.150000 ;
        RECT 1151.000000 493.850000 1156.000000 494.150000 ;
        RECT 1151.000000 497.850000 1156.000000 498.150000 ;
        RECT 1151.000000 505.850000 1156.000000 506.150000 ;
        RECT 1151.000000 501.850000 1156.000000 502.150000 ;
        RECT 1151.000000 509.850000 1156.000000 510.150000 ;
        RECT 1151.000000 513.850000 1156.000000 514.150000 ;
        RECT 1151.000000 517.850000 1156.000000 518.150000 ;
        RECT 1151.000000 521.850000 1156.000000 522.150000 ;
        RECT 1151.000000 525.850000 1156.000000 526.150000 ;
        RECT 1151.000000 533.850000 1156.000000 534.150000 ;
        RECT 1151.000000 529.850000 1156.000000 530.150000 ;
        RECT 1151.000000 545.850000 1156.000000 546.150000 ;
        RECT 1151.000000 537.850000 1156.000000 538.150000 ;
        RECT 1151.000000 541.850000 1156.000000 542.150000 ;
        RECT 1151.000000 553.850000 1156.000000 554.150000 ;
        RECT 1151.000000 549.850000 1156.000000 550.150000 ;
        RECT 1151.000000 561.850000 1156.000000 562.150000 ;
        RECT 1151.000000 557.850000 1156.000000 558.150000 ;
        RECT 1151.000000 565.850000 1156.000000 566.150000 ;
        RECT 1151.000000 569.850000 1156.000000 570.150000 ;
        RECT 1151.000000 573.850000 1156.000000 574.150000 ;
        RECT 1151.000000 577.850000 1156.000000 578.150000 ;
        RECT 1151.000000 581.850000 1156.000000 582.150000 ;
        RECT 1151.000000 589.850000 1156.000000 590.150000 ;
        RECT 1151.000000 585.850000 1156.000000 586.150000 ;
        RECT 1151.000000 593.850000 1156.000000 594.150000 ;
        RECT 1151.000000 597.850000 1156.000000 598.150000 ;
        RECT 1151.000000 601.850000 1156.000000 602.150000 ;
        RECT 1151.000000 609.850000 1156.000000 610.150000 ;
        RECT 1151.000000 605.850000 1156.000000 606.150000 ;
        RECT 1151.000000 613.850000 1156.000000 614.150000 ;
        RECT 1151.000000 617.850000 1156.000000 618.150000 ;
        RECT 1151.000000 621.850000 1156.000000 622.150000 ;
        RECT 1151.000000 625.850000 1156.000000 626.150000 ;
        RECT 1151.000000 629.850000 1156.000000 630.150000 ;
        RECT 1151.000000 637.850000 1156.000000 638.150000 ;
        RECT 1151.000000 633.850000 1156.000000 634.150000 ;
        RECT 601.000000 657.850000 606.000000 658.150000 ;
        RECT 601.000000 673.850000 606.000000 674.150000 ;
        RECT 601.000000 669.850000 606.000000 670.150000 ;
        RECT 601.000000 665.850000 606.000000 666.150000 ;
        RECT 601.000000 661.850000 606.000000 662.150000 ;
        RECT 651.000000 657.850000 656.000000 658.150000 ;
        RECT 651.000000 665.850000 656.000000 666.150000 ;
        RECT 651.000000 661.850000 656.000000 662.150000 ;
        RECT 651.000000 673.850000 656.000000 674.150000 ;
        RECT 651.000000 669.850000 656.000000 670.150000 ;
        RECT 601.000000 677.850000 606.000000 678.150000 ;
        RECT 601.000000 681.850000 606.000000 682.150000 ;
        RECT 651.000000 677.850000 656.000000 678.150000 ;
        RECT 651.000000 681.850000 656.000000 682.150000 ;
        RECT 1151.000000 657.850000 1156.000000 658.150000 ;
        RECT 1151.000000 641.850000 1156.000000 642.150000 ;
        RECT 1151.000000 645.850000 1156.000000 646.150000 ;
        RECT 1151.000000 649.850000 1156.000000 650.150000 ;
        RECT 1151.000000 653.850000 1156.000000 654.150000 ;
        RECT 1151.000000 665.850000 1156.000000 666.150000 ;
        RECT 1151.000000 661.850000 1156.000000 662.150000 ;
        RECT 1151.000000 669.850000 1156.000000 670.150000 ;
        RECT 1151.000000 673.850000 1156.000000 674.150000 ;
        RECT 1151.000000 681.850000 1156.000000 682.150000 ;
        RECT 1151.000000 677.850000 1156.000000 678.150000 ;
      LAYER M3 ;
        RECT 4.000000 5.850000 14.000000 6.150000 ;
        RECT 51.000000 5.850000 56.000000 6.150000 ;
        RECT 51.000000 1.850000 56.000000 2.150000 ;
        RECT 101.000000 1.850000 106.000000 2.150000 ;
        RECT 101.000000 5.850000 106.000000 6.150000 ;
        RECT 151.000000 1.850000 156.000000 2.150000 ;
        RECT 151.000000 5.850000 156.000000 6.150000 ;
        RECT 201.000000 1.850000 206.000000 2.150000 ;
        RECT 201.000000 5.850000 206.000000 6.150000 ;
        RECT 251.000000 1.850000 256.000000 2.150000 ;
        RECT 251.000000 5.850000 256.000000 6.150000 ;
        RECT 301.000000 1.850000 306.000000 2.150000 ;
        RECT 301.000000 5.850000 306.000000 6.150000 ;
        RECT 351.000000 1.850000 356.000000 2.150000 ;
        RECT 351.000000 5.850000 356.000000 6.150000 ;
        RECT 401.000000 1.850000 406.000000 2.150000 ;
        RECT 401.000000 5.850000 406.000000 6.150000 ;
        RECT 451.000000 1.850000 456.000000 2.150000 ;
        RECT 451.000000 5.850000 456.000000 6.150000 ;
        RECT 501.000000 1.850000 506.000000 2.150000 ;
        RECT 501.000000 5.850000 506.000000 6.150000 ;
        RECT 551.000000 1.850000 556.000000 2.150000 ;
        RECT 551.000000 5.850000 556.000000 6.150000 ;
        RECT 4.000000 265.850000 14.000000 266.150000 ;
        RECT 4.000000 261.850000 14.000000 262.150000 ;
        RECT 51.000000 265.850000 56.000000 266.150000 ;
        RECT 51.000000 261.850000 56.000000 262.150000 ;
        RECT 101.000000 265.850000 106.000000 266.150000 ;
        RECT 101.000000 261.850000 106.000000 262.150000 ;
        RECT 51.000000 305.850000 56.000000 306.150000 ;
        RECT 4.000000 305.850000 14.000000 306.150000 ;
        RECT 4.000000 285.850000 14.000000 286.150000 ;
        RECT 4.000000 281.850000 14.000000 282.150000 ;
        RECT 4.000000 269.850000 14.000000 270.150000 ;
        RECT 4.000000 273.850000 14.000000 274.150000 ;
        RECT 4.000000 277.850000 14.000000 278.150000 ;
        RECT 4.000000 289.850000 14.000000 290.150000 ;
        RECT 4.000000 293.850000 14.000000 294.150000 ;
        RECT 4.000000 297.850000 14.000000 298.150000 ;
        RECT 4.000000 301.850000 14.000000 302.150000 ;
        RECT 51.000000 269.850000 56.000000 270.150000 ;
        RECT 51.000000 273.850000 56.000000 274.150000 ;
        RECT 51.000000 277.850000 56.000000 278.150000 ;
        RECT 51.000000 281.850000 56.000000 282.150000 ;
        RECT 51.000000 285.850000 56.000000 286.150000 ;
        RECT 51.000000 301.850000 56.000000 302.150000 ;
        RECT 51.000000 297.850000 56.000000 298.150000 ;
        RECT 51.000000 293.850000 56.000000 294.150000 ;
        RECT 51.000000 289.850000 56.000000 290.150000 ;
        RECT 4.000000 321.850000 14.000000 322.150000 ;
        RECT 4.000000 309.850000 14.000000 310.150000 ;
        RECT 4.000000 313.850000 14.000000 314.150000 ;
        RECT 4.000000 317.850000 14.000000 318.150000 ;
        RECT 4.000000 325.850000 14.000000 326.150000 ;
        RECT 4.000000 329.850000 14.000000 330.150000 ;
        RECT 4.000000 333.850000 14.000000 334.150000 ;
        RECT 4.000000 337.850000 14.000000 338.150000 ;
        RECT 4.000000 341.850000 14.000000 342.150000 ;
        RECT 51.000000 313.850000 56.000000 314.150000 ;
        RECT 51.000000 309.850000 56.000000 310.150000 ;
        RECT 51.000000 317.850000 56.000000 318.150000 ;
        RECT 51.000000 321.850000 56.000000 322.150000 ;
        RECT 51.000000 341.850000 56.000000 342.150000 ;
        RECT 51.000000 337.850000 56.000000 338.150000 ;
        RECT 51.000000 333.850000 56.000000 334.150000 ;
        RECT 51.000000 329.850000 56.000000 330.150000 ;
        RECT 51.000000 325.850000 56.000000 326.150000 ;
        RECT 101.000000 305.850000 106.000000 306.150000 ;
        RECT 101.000000 269.850000 106.000000 270.150000 ;
        RECT 101.000000 273.850000 106.000000 274.150000 ;
        RECT 101.000000 277.850000 106.000000 278.150000 ;
        RECT 101.000000 281.850000 106.000000 282.150000 ;
        RECT 101.000000 285.850000 106.000000 286.150000 ;
        RECT 101.000000 301.850000 106.000000 302.150000 ;
        RECT 101.000000 297.850000 106.000000 298.150000 ;
        RECT 101.000000 293.850000 106.000000 294.150000 ;
        RECT 101.000000 289.850000 106.000000 290.150000 ;
        RECT 101.000000 321.850000 106.000000 322.150000 ;
        RECT 101.000000 317.850000 106.000000 318.150000 ;
        RECT 101.000000 313.850000 106.000000 314.150000 ;
        RECT 101.000000 309.850000 106.000000 310.150000 ;
        RECT 101.000000 325.850000 106.000000 326.150000 ;
        RECT 101.000000 329.850000 106.000000 330.150000 ;
        RECT 101.000000 333.850000 106.000000 334.150000 ;
        RECT 101.000000 337.850000 106.000000 338.150000 ;
        RECT 101.000000 341.850000 106.000000 342.150000 ;
        RECT 151.000000 261.850000 156.000000 262.150000 ;
        RECT 151.000000 265.850000 156.000000 266.150000 ;
        RECT 201.000000 265.850000 206.000000 266.150000 ;
        RECT 201.000000 261.850000 206.000000 262.150000 ;
        RECT 251.000000 265.850000 256.000000 266.150000 ;
        RECT 251.000000 261.850000 256.000000 262.150000 ;
        RECT 201.000000 305.850000 206.000000 306.150000 ;
        RECT 151.000000 305.850000 156.000000 306.150000 ;
        RECT 151.000000 277.850000 156.000000 278.150000 ;
        RECT 151.000000 273.850000 156.000000 274.150000 ;
        RECT 151.000000 269.850000 156.000000 270.150000 ;
        RECT 151.000000 281.850000 156.000000 282.150000 ;
        RECT 151.000000 285.850000 156.000000 286.150000 ;
        RECT 151.000000 289.850000 156.000000 290.150000 ;
        RECT 151.000000 293.850000 156.000000 294.150000 ;
        RECT 151.000000 297.850000 156.000000 298.150000 ;
        RECT 151.000000 301.850000 156.000000 302.150000 ;
        RECT 201.000000 269.850000 206.000000 270.150000 ;
        RECT 201.000000 273.850000 206.000000 274.150000 ;
        RECT 201.000000 277.850000 206.000000 278.150000 ;
        RECT 201.000000 281.850000 206.000000 282.150000 ;
        RECT 201.000000 285.850000 206.000000 286.150000 ;
        RECT 201.000000 301.850000 206.000000 302.150000 ;
        RECT 201.000000 297.850000 206.000000 298.150000 ;
        RECT 201.000000 293.850000 206.000000 294.150000 ;
        RECT 201.000000 289.850000 206.000000 290.150000 ;
        RECT 151.000000 313.850000 156.000000 314.150000 ;
        RECT 151.000000 309.850000 156.000000 310.150000 ;
        RECT 151.000000 321.850000 156.000000 322.150000 ;
        RECT 151.000000 317.850000 156.000000 318.150000 ;
        RECT 151.000000 329.850000 156.000000 330.150000 ;
        RECT 151.000000 325.850000 156.000000 326.150000 ;
        RECT 151.000000 333.850000 156.000000 334.150000 ;
        RECT 151.000000 337.850000 156.000000 338.150000 ;
        RECT 151.000000 341.850000 156.000000 342.150000 ;
        RECT 201.000000 313.850000 206.000000 314.150000 ;
        RECT 201.000000 309.850000 206.000000 310.150000 ;
        RECT 201.000000 317.850000 206.000000 318.150000 ;
        RECT 201.000000 321.850000 206.000000 322.150000 ;
        RECT 201.000000 341.850000 206.000000 342.150000 ;
        RECT 201.000000 337.850000 206.000000 338.150000 ;
        RECT 201.000000 333.850000 206.000000 334.150000 ;
        RECT 201.000000 329.850000 206.000000 330.150000 ;
        RECT 201.000000 325.850000 206.000000 326.150000 ;
        RECT 251.000000 305.850000 256.000000 306.150000 ;
        RECT 251.000000 269.850000 256.000000 270.150000 ;
        RECT 251.000000 273.850000 256.000000 274.150000 ;
        RECT 251.000000 277.850000 256.000000 278.150000 ;
        RECT 251.000000 281.850000 256.000000 282.150000 ;
        RECT 251.000000 285.850000 256.000000 286.150000 ;
        RECT 251.000000 293.850000 256.000000 294.150000 ;
        RECT 251.000000 289.850000 256.000000 290.150000 ;
        RECT 251.000000 301.850000 256.000000 302.150000 ;
        RECT 251.000000 297.850000 256.000000 298.150000 ;
        RECT 251.000000 321.850000 256.000000 322.150000 ;
        RECT 251.000000 317.850000 256.000000 318.150000 ;
        RECT 251.000000 313.850000 256.000000 314.150000 ;
        RECT 251.000000 309.850000 256.000000 310.150000 ;
        RECT 251.000000 325.850000 256.000000 326.150000 ;
        RECT 251.000000 329.850000 256.000000 330.150000 ;
        RECT 251.000000 337.850000 256.000000 338.150000 ;
        RECT 251.000000 333.850000 256.000000 334.150000 ;
        RECT 251.000000 341.850000 256.000000 342.150000 ;
        RECT 301.000000 265.850000 306.000000 266.150000 ;
        RECT 301.000000 261.850000 306.000000 262.150000 ;
        RECT 351.000000 265.850000 356.000000 266.150000 ;
        RECT 351.000000 261.850000 356.000000 262.150000 ;
        RECT 401.000000 261.850000 406.000000 262.150000 ;
        RECT 401.000000 265.850000 406.000000 266.150000 ;
        RECT 351.000000 305.850000 356.000000 306.150000 ;
        RECT 301.000000 305.850000 306.000000 306.150000 ;
        RECT 301.000000 277.850000 306.000000 278.150000 ;
        RECT 301.000000 269.850000 306.000000 270.150000 ;
        RECT 301.000000 273.850000 306.000000 274.150000 ;
        RECT 301.000000 281.850000 306.000000 282.150000 ;
        RECT 301.000000 285.850000 306.000000 286.150000 ;
        RECT 301.000000 293.850000 306.000000 294.150000 ;
        RECT 301.000000 289.850000 306.000000 290.150000 ;
        RECT 301.000000 301.850000 306.000000 302.150000 ;
        RECT 301.000000 297.850000 306.000000 298.150000 ;
        RECT 351.000000 269.850000 356.000000 270.150000 ;
        RECT 351.000000 273.850000 356.000000 274.150000 ;
        RECT 351.000000 277.850000 356.000000 278.150000 ;
        RECT 351.000000 281.850000 356.000000 282.150000 ;
        RECT 351.000000 285.850000 356.000000 286.150000 ;
        RECT 351.000000 301.850000 356.000000 302.150000 ;
        RECT 351.000000 297.850000 356.000000 298.150000 ;
        RECT 351.000000 293.850000 356.000000 294.150000 ;
        RECT 351.000000 289.850000 356.000000 290.150000 ;
        RECT 301.000000 313.850000 306.000000 314.150000 ;
        RECT 301.000000 309.850000 306.000000 310.150000 ;
        RECT 301.000000 317.850000 306.000000 318.150000 ;
        RECT 301.000000 321.850000 306.000000 322.150000 ;
        RECT 301.000000 329.850000 306.000000 330.150000 ;
        RECT 301.000000 325.850000 306.000000 326.150000 ;
        RECT 301.000000 341.850000 306.000000 342.150000 ;
        RECT 301.000000 337.850000 306.000000 338.150000 ;
        RECT 301.000000 333.850000 306.000000 334.150000 ;
        RECT 351.000000 313.850000 356.000000 314.150000 ;
        RECT 351.000000 309.850000 356.000000 310.150000 ;
        RECT 351.000000 317.850000 356.000000 318.150000 ;
        RECT 351.000000 321.850000 356.000000 322.150000 ;
        RECT 351.000000 341.850000 356.000000 342.150000 ;
        RECT 351.000000 337.850000 356.000000 338.150000 ;
        RECT 351.000000 333.850000 356.000000 334.150000 ;
        RECT 351.000000 329.850000 356.000000 330.150000 ;
        RECT 351.000000 325.850000 356.000000 326.150000 ;
        RECT 401.000000 305.850000 406.000000 306.150000 ;
        RECT 401.000000 277.850000 406.000000 278.150000 ;
        RECT 401.000000 269.850000 406.000000 270.150000 ;
        RECT 401.000000 273.850000 406.000000 274.150000 ;
        RECT 401.000000 281.850000 406.000000 282.150000 ;
        RECT 401.000000 285.850000 406.000000 286.150000 ;
        RECT 401.000000 301.850000 406.000000 302.150000 ;
        RECT 401.000000 297.850000 406.000000 298.150000 ;
        RECT 401.000000 293.850000 406.000000 294.150000 ;
        RECT 401.000000 289.850000 406.000000 290.150000 ;
        RECT 401.000000 313.850000 406.000000 314.150000 ;
        RECT 401.000000 309.850000 406.000000 310.150000 ;
        RECT 401.000000 317.850000 406.000000 318.150000 ;
        RECT 401.000000 321.850000 406.000000 322.150000 ;
        RECT 401.000000 329.850000 406.000000 330.150000 ;
        RECT 401.000000 325.850000 406.000000 326.150000 ;
        RECT 401.000000 333.850000 406.000000 334.150000 ;
        RECT 401.000000 337.850000 406.000000 338.150000 ;
        RECT 401.000000 341.850000 406.000000 342.150000 ;
        RECT 451.000000 265.850000 456.000000 266.150000 ;
        RECT 451.000000 261.850000 456.000000 262.150000 ;
        RECT 501.000000 261.850000 506.000000 262.150000 ;
        RECT 501.000000 265.850000 506.000000 266.150000 ;
        RECT 551.000000 265.850000 556.000000 266.150000 ;
        RECT 551.000000 261.850000 556.000000 262.150000 ;
        RECT 501.000000 305.850000 506.000000 306.150000 ;
        RECT 451.000000 277.850000 456.000000 278.150000 ;
        RECT 451.000000 273.850000 456.000000 274.150000 ;
        RECT 451.000000 269.850000 456.000000 270.150000 ;
        RECT 451.000000 285.850000 456.000000 286.150000 ;
        RECT 451.000000 281.850000 456.000000 282.150000 ;
        RECT 451.000000 293.850000 456.000000 294.150000 ;
        RECT 451.000000 289.850000 456.000000 290.150000 ;
        RECT 451.000000 297.850000 456.000000 298.150000 ;
        RECT 501.000000 277.850000 506.000000 278.150000 ;
        RECT 501.000000 269.850000 506.000000 270.150000 ;
        RECT 501.000000 273.850000 506.000000 274.150000 ;
        RECT 501.000000 281.850000 506.000000 282.150000 ;
        RECT 501.000000 285.850000 506.000000 286.150000 ;
        RECT 501.000000 289.850000 506.000000 290.150000 ;
        RECT 501.000000 293.850000 506.000000 294.150000 ;
        RECT 501.000000 297.850000 506.000000 298.150000 ;
        RECT 501.000000 301.850000 506.000000 302.150000 ;
        RECT 451.000000 316.105000 456.000000 317.105000 ;
        RECT 451.000000 321.850000 456.000000 322.150000 ;
        RECT 451.000000 333.850000 456.000000 334.150000 ;
        RECT 451.000000 329.850000 456.000000 330.150000 ;
        RECT 451.000000 325.850000 456.000000 326.150000 ;
        RECT 451.000000 337.850000 456.000000 338.150000 ;
        RECT 451.000000 341.850000 456.000000 342.150000 ;
        RECT 501.000000 313.850000 506.000000 314.150000 ;
        RECT 501.000000 309.850000 506.000000 310.150000 ;
        RECT 501.000000 317.850000 506.000000 318.150000 ;
        RECT 501.000000 321.850000 506.000000 322.150000 ;
        RECT 501.000000 329.850000 506.000000 330.150000 ;
        RECT 501.000000 325.850000 506.000000 326.150000 ;
        RECT 501.000000 333.850000 506.000000 334.150000 ;
        RECT 501.000000 337.850000 506.000000 338.150000 ;
        RECT 501.000000 341.850000 506.000000 342.150000 ;
        RECT 551.000000 305.850000 556.000000 306.150000 ;
        RECT 551.000000 285.850000 556.000000 286.150000 ;
        RECT 551.000000 281.850000 556.000000 282.150000 ;
        RECT 551.000000 277.850000 556.000000 278.150000 ;
        RECT 551.000000 273.850000 556.000000 274.150000 ;
        RECT 551.000000 269.850000 556.000000 270.150000 ;
        RECT 551.000000 301.850000 556.000000 302.150000 ;
        RECT 551.000000 297.850000 556.000000 298.150000 ;
        RECT 551.000000 293.850000 556.000000 294.150000 ;
        RECT 551.000000 289.850000 556.000000 290.150000 ;
        RECT 551.000000 309.850000 556.000000 310.150000 ;
        RECT 551.000000 313.850000 556.000000 314.150000 ;
        RECT 551.000000 317.850000 556.000000 318.150000 ;
        RECT 551.000000 321.850000 556.000000 322.150000 ;
        RECT 551.000000 325.850000 556.000000 326.150000 ;
        RECT 551.000000 329.850000 556.000000 330.150000 ;
        RECT 551.000000 333.850000 556.000000 334.150000 ;
        RECT 551.000000 337.850000 556.000000 338.150000 ;
        RECT 551.000000 341.850000 556.000000 342.150000 ;
        RECT 601.000000 1.850000 606.000000 2.150000 ;
        RECT 601.000000 5.850000 606.000000 6.150000 ;
        RECT 651.000000 1.850000 656.000000 2.150000 ;
        RECT 651.000000 5.850000 656.000000 6.150000 ;
        RECT 701.000000 1.850000 706.000000 2.150000 ;
        RECT 701.000000 5.850000 706.000000 6.150000 ;
        RECT 751.000000 1.850000 756.000000 2.150000 ;
        RECT 751.000000 5.850000 756.000000 6.150000 ;
        RECT 801.000000 1.850000 806.000000 2.150000 ;
        RECT 801.000000 5.850000 806.000000 6.150000 ;
        RECT 851.000000 1.850000 856.000000 2.150000 ;
        RECT 851.000000 5.850000 856.000000 6.150000 ;
        RECT 901.000000 1.850000 906.000000 2.150000 ;
        RECT 901.000000 5.850000 906.000000 6.150000 ;
        RECT 951.000000 1.850000 956.000000 2.150000 ;
        RECT 951.000000 5.850000 956.000000 6.150000 ;
        RECT 1001.000000 1.850000 1006.000000 2.150000 ;
        RECT 1001.000000 5.850000 1006.000000 6.150000 ;
        RECT 1051.000000 1.850000 1056.000000 2.150000 ;
        RECT 1051.000000 5.850000 1056.000000 6.150000 ;
        RECT 1101.000000 1.850000 1106.000000 2.150000 ;
        RECT 1101.000000 5.850000 1106.000000 6.150000 ;
        RECT 1151.000000 5.850000 1156.000000 6.150000 ;
        RECT 1172.000000 5.850000 1182.000000 6.150000 ;
        RECT 1151.000000 1.850000 1156.000000 2.150000 ;
        RECT 1172.000000 17.850000 1182.000000 18.150000 ;
        RECT 1172.000000 13.850000 1182.000000 14.150000 ;
        RECT 1172.000000 9.850000 1182.000000 10.150000 ;
        RECT 1172.000000 21.850000 1182.000000 22.150000 ;
        RECT 1172.000000 25.850000 1182.000000 26.150000 ;
        RECT 1172.000000 33.850000 1182.000000 34.150000 ;
        RECT 1172.000000 29.850000 1182.000000 30.150000 ;
        RECT 1172.000000 41.850000 1182.000000 42.150000 ;
        RECT 1172.000000 37.850000 1182.000000 38.150000 ;
        RECT 1172.000000 45.850000 1182.000000 46.150000 ;
        RECT 601.000000 261.850000 606.000000 262.150000 ;
        RECT 601.000000 265.850000 606.000000 266.150000 ;
        RECT 651.000000 261.850000 656.000000 262.150000 ;
        RECT 651.000000 265.850000 656.000000 266.150000 ;
        RECT 701.000000 265.850000 706.000000 266.150000 ;
        RECT 701.000000 261.850000 706.000000 262.150000 ;
        RECT 601.000000 305.850000 606.000000 306.150000 ;
        RECT 651.000000 305.850000 656.000000 306.150000 ;
        RECT 601.000000 277.850000 606.000000 278.150000 ;
        RECT 601.000000 269.850000 606.000000 270.150000 ;
        RECT 601.000000 273.850000 606.000000 274.150000 ;
        RECT 601.000000 281.850000 606.000000 282.150000 ;
        RECT 601.000000 285.850000 606.000000 286.150000 ;
        RECT 601.000000 289.850000 606.000000 290.150000 ;
        RECT 601.000000 293.850000 606.000000 294.150000 ;
        RECT 601.000000 297.850000 606.000000 298.150000 ;
        RECT 601.000000 301.850000 606.000000 302.150000 ;
        RECT 651.000000 277.850000 656.000000 278.150000 ;
        RECT 651.000000 273.850000 656.000000 274.150000 ;
        RECT 651.000000 269.850000 656.000000 270.150000 ;
        RECT 651.000000 281.850000 656.000000 282.150000 ;
        RECT 651.000000 285.850000 656.000000 286.150000 ;
        RECT 651.000000 289.850000 656.000000 290.150000 ;
        RECT 651.000000 293.850000 656.000000 294.150000 ;
        RECT 651.000000 301.850000 656.000000 302.150000 ;
        RECT 651.000000 297.850000 656.000000 298.150000 ;
        RECT 601.000000 321.850000 606.000000 322.150000 ;
        RECT 601.000000 317.850000 606.000000 318.150000 ;
        RECT 601.000000 309.850000 606.000000 310.150000 ;
        RECT 601.000000 313.850000 606.000000 314.150000 ;
        RECT 601.000000 325.850000 606.000000 326.150000 ;
        RECT 601.000000 329.850000 606.000000 330.150000 ;
        RECT 601.000000 333.850000 606.000000 334.150000 ;
        RECT 601.000000 337.850000 606.000000 338.150000 ;
        RECT 601.000000 341.850000 606.000000 342.150000 ;
        RECT 651.000000 313.850000 656.000000 314.150000 ;
        RECT 651.000000 309.850000 656.000000 310.150000 ;
        RECT 651.000000 321.850000 656.000000 322.150000 ;
        RECT 651.000000 317.850000 656.000000 318.150000 ;
        RECT 651.000000 329.850000 656.000000 330.150000 ;
        RECT 651.000000 325.850000 656.000000 326.150000 ;
        RECT 651.000000 333.850000 656.000000 334.150000 ;
        RECT 651.000000 337.850000 656.000000 338.150000 ;
        RECT 651.000000 341.850000 656.000000 342.150000 ;
        RECT 701.000000 305.850000 706.000000 306.150000 ;
        RECT 701.000000 285.850000 706.000000 286.150000 ;
        RECT 701.000000 281.850000 706.000000 282.150000 ;
        RECT 701.000000 277.850000 706.000000 278.150000 ;
        RECT 701.000000 273.850000 706.000000 274.150000 ;
        RECT 701.000000 269.850000 706.000000 270.150000 ;
        RECT 701.000000 301.850000 706.000000 302.150000 ;
        RECT 701.000000 297.850000 706.000000 298.150000 ;
        RECT 701.000000 293.850000 706.000000 294.150000 ;
        RECT 701.000000 289.850000 706.000000 290.150000 ;
        RECT 701.000000 309.850000 706.000000 310.150000 ;
        RECT 701.000000 313.850000 706.000000 314.150000 ;
        RECT 701.000000 317.850000 706.000000 318.150000 ;
        RECT 701.000000 321.850000 706.000000 322.150000 ;
        RECT 701.000000 325.850000 706.000000 326.150000 ;
        RECT 701.000000 329.850000 706.000000 330.150000 ;
        RECT 701.000000 333.850000 706.000000 334.150000 ;
        RECT 701.000000 337.850000 706.000000 338.150000 ;
        RECT 701.000000 341.850000 706.000000 342.150000 ;
        RECT 751.000000 261.850000 756.000000 262.150000 ;
        RECT 751.000000 265.850000 756.000000 266.150000 ;
        RECT 801.000000 261.850000 806.000000 262.150000 ;
        RECT 801.000000 265.850000 806.000000 266.150000 ;
        RECT 851.000000 265.850000 856.000000 266.150000 ;
        RECT 851.000000 261.850000 856.000000 262.150000 ;
        RECT 801.000000 305.850000 806.000000 306.150000 ;
        RECT 751.000000 305.850000 756.000000 306.150000 ;
        RECT 751.000000 285.850000 756.000000 286.150000 ;
        RECT 751.000000 281.850000 756.000000 282.150000 ;
        RECT 751.000000 269.850000 756.000000 270.150000 ;
        RECT 751.000000 273.850000 756.000000 274.150000 ;
        RECT 751.000000 277.850000 756.000000 278.150000 ;
        RECT 751.000000 289.850000 756.000000 290.150000 ;
        RECT 751.000000 293.850000 756.000000 294.150000 ;
        RECT 751.000000 297.850000 756.000000 298.150000 ;
        RECT 751.000000 301.850000 756.000000 302.150000 ;
        RECT 801.000000 277.850000 806.000000 278.150000 ;
        RECT 801.000000 269.850000 806.000000 270.150000 ;
        RECT 801.000000 273.850000 806.000000 274.150000 ;
        RECT 801.000000 281.850000 806.000000 282.150000 ;
        RECT 801.000000 285.850000 806.000000 286.150000 ;
        RECT 801.000000 289.850000 806.000000 290.150000 ;
        RECT 801.000000 293.850000 806.000000 294.150000 ;
        RECT 801.000000 301.850000 806.000000 302.150000 ;
        RECT 801.000000 297.850000 806.000000 298.150000 ;
        RECT 751.000000 321.850000 756.000000 322.150000 ;
        RECT 751.000000 309.850000 756.000000 310.150000 ;
        RECT 751.000000 313.850000 756.000000 314.150000 ;
        RECT 751.000000 317.850000 756.000000 318.150000 ;
        RECT 751.000000 325.850000 756.000000 326.150000 ;
        RECT 751.000000 329.850000 756.000000 330.150000 ;
        RECT 751.000000 333.850000 756.000000 334.150000 ;
        RECT 751.000000 337.850000 756.000000 338.150000 ;
        RECT 751.000000 341.850000 756.000000 342.150000 ;
        RECT 801.000000 313.850000 806.000000 314.150000 ;
        RECT 801.000000 309.850000 806.000000 310.150000 ;
        RECT 801.000000 321.850000 806.000000 322.150000 ;
        RECT 801.000000 317.850000 806.000000 318.150000 ;
        RECT 801.000000 329.850000 806.000000 330.150000 ;
        RECT 801.000000 325.850000 806.000000 326.150000 ;
        RECT 801.000000 333.850000 806.000000 334.150000 ;
        RECT 801.000000 337.850000 806.000000 338.150000 ;
        RECT 801.000000 341.850000 806.000000 342.150000 ;
        RECT 851.000000 305.850000 856.000000 306.150000 ;
        RECT 851.000000 285.850000 856.000000 286.150000 ;
        RECT 851.000000 281.850000 856.000000 282.150000 ;
        RECT 851.000000 277.850000 856.000000 278.150000 ;
        RECT 851.000000 273.850000 856.000000 274.150000 ;
        RECT 851.000000 269.850000 856.000000 270.150000 ;
        RECT 851.000000 301.850000 856.000000 302.150000 ;
        RECT 851.000000 297.850000 856.000000 298.150000 ;
        RECT 851.000000 293.850000 856.000000 294.150000 ;
        RECT 851.000000 289.850000 856.000000 290.150000 ;
        RECT 851.000000 309.850000 856.000000 310.150000 ;
        RECT 851.000000 313.850000 856.000000 314.150000 ;
        RECT 851.000000 317.850000 856.000000 318.150000 ;
        RECT 851.000000 321.850000 856.000000 322.150000 ;
        RECT 851.000000 325.850000 856.000000 326.150000 ;
        RECT 851.000000 329.850000 856.000000 330.150000 ;
        RECT 851.000000 333.850000 856.000000 334.150000 ;
        RECT 851.000000 337.850000 856.000000 338.150000 ;
        RECT 851.000000 341.850000 856.000000 342.150000 ;
        RECT 1172.000000 61.850000 1182.000000 62.150000 ;
        RECT 1172.000000 57.850000 1182.000000 58.150000 ;
        RECT 1172.000000 53.850000 1182.000000 54.150000 ;
        RECT 1172.000000 49.850000 1182.000000 50.150000 ;
        RECT 1172.000000 73.850000 1182.000000 74.150000 ;
        RECT 1172.000000 69.850000 1182.000000 70.150000 ;
        RECT 1172.000000 65.850000 1182.000000 66.150000 ;
        RECT 1172.000000 77.850000 1182.000000 78.150000 ;
        RECT 1172.000000 81.850000 1182.000000 82.150000 ;
        RECT 1172.000000 101.850000 1182.000000 102.150000 ;
        RECT 1172.000000 85.850000 1182.000000 86.150000 ;
        RECT 1172.000000 89.850000 1182.000000 90.150000 ;
        RECT 1172.000000 93.850000 1182.000000 94.150000 ;
        RECT 1172.000000 97.850000 1182.000000 98.150000 ;
        RECT 1172.000000 117.850000 1182.000000 118.150000 ;
        RECT 1172.000000 113.850000 1182.000000 114.150000 ;
        RECT 1172.000000 105.850000 1182.000000 106.150000 ;
        RECT 1172.000000 109.850000 1182.000000 110.150000 ;
        RECT 1151.000000 133.850000 1156.000000 134.150000 ;
        RECT 1172.000000 129.850000 1182.000000 130.150000 ;
        RECT 1172.000000 125.850000 1182.000000 126.150000 ;
        RECT 1172.000000 121.850000 1182.000000 122.150000 ;
        RECT 1172.000000 133.850000 1182.000000 134.150000 ;
        RECT 1172.000000 137.850000 1182.000000 138.150000 ;
        RECT 1172.000000 141.850000 1182.000000 142.150000 ;
        RECT 1172.000000 145.850000 1182.000000 146.150000 ;
        RECT 1172.000000 149.850000 1182.000000 150.150000 ;
        RECT 1172.000000 153.850000 1182.000000 154.150000 ;
        RECT 1172.000000 165.850000 1182.000000 166.150000 ;
        RECT 1172.000000 161.850000 1182.000000 162.150000 ;
        RECT 1172.000000 157.850000 1182.000000 158.150000 ;
        RECT 1172.000000 169.850000 1182.000000 170.150000 ;
        RECT 1172.000000 173.850000 1182.000000 174.150000 ;
        RECT 1172.000000 177.850000 1182.000000 178.150000 ;
        RECT 1172.000000 181.850000 1182.000000 182.150000 ;
        RECT 1172.000000 185.850000 1182.000000 186.150000 ;
        RECT 1172.000000 189.850000 1182.000000 190.150000 ;
        RECT 1172.000000 193.850000 1182.000000 194.150000 ;
        RECT 901.000000 261.850000 906.000000 262.150000 ;
        RECT 901.000000 265.850000 906.000000 266.150000 ;
        RECT 951.000000 265.850000 956.000000 266.150000 ;
        RECT 951.000000 261.850000 956.000000 262.150000 ;
        RECT 1001.000000 261.850000 1006.000000 262.150000 ;
        RECT 1001.000000 265.850000 1006.000000 266.150000 ;
        RECT 951.000000 305.850000 956.000000 306.150000 ;
        RECT 901.000000 305.850000 906.000000 306.150000 ;
        RECT 901.000000 285.850000 906.000000 286.150000 ;
        RECT 901.000000 281.850000 906.000000 282.150000 ;
        RECT 901.000000 269.850000 906.000000 270.150000 ;
        RECT 901.000000 273.850000 906.000000 274.150000 ;
        RECT 901.000000 277.850000 906.000000 278.150000 ;
        RECT 901.000000 289.850000 906.000000 290.150000 ;
        RECT 901.000000 293.850000 906.000000 294.150000 ;
        RECT 901.000000 297.850000 906.000000 298.150000 ;
        RECT 901.000000 301.850000 906.000000 302.150000 ;
        RECT 951.000000 269.850000 956.000000 270.150000 ;
        RECT 951.000000 273.850000 956.000000 274.150000 ;
        RECT 951.000000 277.850000 956.000000 278.150000 ;
        RECT 951.000000 281.850000 956.000000 282.150000 ;
        RECT 951.000000 285.850000 956.000000 286.150000 ;
        RECT 951.000000 301.850000 956.000000 302.150000 ;
        RECT 951.000000 297.850000 956.000000 298.150000 ;
        RECT 951.000000 293.850000 956.000000 294.150000 ;
        RECT 951.000000 289.850000 956.000000 290.150000 ;
        RECT 901.000000 321.850000 906.000000 322.150000 ;
        RECT 901.000000 309.850000 906.000000 310.150000 ;
        RECT 901.000000 313.850000 906.000000 314.150000 ;
        RECT 901.000000 317.850000 906.000000 318.150000 ;
        RECT 901.000000 325.850000 906.000000 326.150000 ;
        RECT 901.000000 329.850000 906.000000 330.150000 ;
        RECT 901.000000 333.850000 906.000000 334.150000 ;
        RECT 901.000000 337.850000 906.000000 338.150000 ;
        RECT 901.000000 341.850000 906.000000 342.150000 ;
        RECT 951.000000 313.850000 956.000000 314.150000 ;
        RECT 951.000000 309.850000 956.000000 310.150000 ;
        RECT 951.000000 317.850000 956.000000 318.150000 ;
        RECT 951.000000 321.850000 956.000000 322.150000 ;
        RECT 951.000000 325.850000 956.000000 326.150000 ;
        RECT 951.000000 329.850000 956.000000 330.150000 ;
        RECT 951.000000 333.850000 956.000000 334.150000 ;
        RECT 951.000000 337.850000 956.000000 338.150000 ;
        RECT 951.000000 341.850000 956.000000 342.150000 ;
        RECT 1001.000000 305.850000 1006.000000 306.150000 ;
        RECT 1001.000000 277.850000 1006.000000 278.150000 ;
        RECT 1001.000000 269.850000 1006.000000 270.150000 ;
        RECT 1001.000000 273.850000 1006.000000 274.150000 ;
        RECT 1001.000000 281.850000 1006.000000 282.150000 ;
        RECT 1001.000000 285.850000 1006.000000 286.150000 ;
        RECT 1001.000000 289.850000 1006.000000 290.150000 ;
        RECT 1001.000000 293.850000 1006.000000 294.150000 ;
        RECT 1001.000000 301.850000 1006.000000 302.150000 ;
        RECT 1001.000000 297.850000 1006.000000 298.150000 ;
        RECT 1001.000000 313.850000 1006.000000 314.150000 ;
        RECT 1001.000000 309.850000 1006.000000 310.150000 ;
        RECT 1001.000000 317.850000 1006.000000 318.150000 ;
        RECT 1001.000000 321.850000 1006.000000 322.150000 ;
        RECT 1001.000000 329.850000 1006.000000 330.150000 ;
        RECT 1001.000000 325.850000 1006.000000 326.150000 ;
        RECT 1001.000000 333.850000 1006.000000 334.150000 ;
        RECT 1001.000000 337.850000 1006.000000 338.150000 ;
        RECT 1001.000000 341.850000 1006.000000 342.150000 ;
        RECT 1051.000000 261.850000 1056.000000 262.150000 ;
        RECT 1051.000000 265.850000 1056.000000 266.150000 ;
        RECT 1101.000000 265.850000 1106.000000 266.150000 ;
        RECT 1101.000000 261.850000 1106.000000 262.150000 ;
        RECT 1172.000000 197.850000 1182.000000 198.150000 ;
        RECT 1172.000000 201.850000 1182.000000 202.150000 ;
        RECT 1172.000000 205.850000 1182.000000 206.150000 ;
        RECT 1172.000000 209.850000 1182.000000 210.150000 ;
        RECT 1172.000000 221.850000 1182.000000 222.150000 ;
        RECT 1172.000000 217.850000 1182.000000 218.150000 ;
        RECT 1172.000000 213.850000 1182.000000 214.150000 ;
        RECT 1172.000000 225.850000 1182.000000 226.150000 ;
        RECT 1172.000000 229.850000 1182.000000 230.150000 ;
        RECT 1172.000000 237.850000 1182.000000 238.150000 ;
        RECT 1172.000000 233.850000 1182.000000 234.150000 ;
        RECT 1172.000000 241.850000 1182.000000 242.150000 ;
        RECT 1172.000000 245.850000 1182.000000 246.150000 ;
        RECT 1172.000000 249.850000 1182.000000 250.150000 ;
        RECT 1151.000000 257.850000 1156.000000 258.150000 ;
        RECT 1151.000000 265.850000 1156.000000 266.150000 ;
        RECT 1151.000000 261.850000 1156.000000 262.150000 ;
        RECT 1172.000000 265.850000 1182.000000 266.150000 ;
        RECT 1172.000000 253.850000 1182.000000 254.150000 ;
        RECT 1172.000000 257.850000 1182.000000 258.150000 ;
        RECT 1172.000000 261.850000 1182.000000 262.150000 ;
        RECT 1101.000000 305.850000 1106.000000 306.150000 ;
        RECT 1051.000000 305.850000 1056.000000 306.150000 ;
        RECT 1051.000000 285.850000 1056.000000 286.150000 ;
        RECT 1051.000000 281.850000 1056.000000 282.150000 ;
        RECT 1051.000000 273.850000 1056.000000 274.150000 ;
        RECT 1051.000000 269.850000 1056.000000 270.150000 ;
        RECT 1051.000000 277.850000 1056.000000 278.150000 ;
        RECT 1051.000000 289.850000 1056.000000 290.150000 ;
        RECT 1051.000000 293.850000 1056.000000 294.150000 ;
        RECT 1051.000000 297.850000 1056.000000 298.150000 ;
        RECT 1051.000000 301.850000 1056.000000 302.150000 ;
        RECT 1101.000000 269.850000 1106.000000 270.150000 ;
        RECT 1101.000000 273.850000 1106.000000 274.150000 ;
        RECT 1101.000000 277.850000 1106.000000 278.150000 ;
        RECT 1101.000000 281.850000 1106.000000 282.150000 ;
        RECT 1101.000000 285.850000 1106.000000 286.150000 ;
        RECT 1101.000000 301.850000 1106.000000 302.150000 ;
        RECT 1101.000000 297.850000 1106.000000 298.150000 ;
        RECT 1101.000000 293.850000 1106.000000 294.150000 ;
        RECT 1101.000000 289.850000 1106.000000 290.150000 ;
        RECT 1051.000000 321.850000 1056.000000 322.150000 ;
        RECT 1051.000000 309.850000 1056.000000 310.150000 ;
        RECT 1051.000000 313.850000 1056.000000 314.150000 ;
        RECT 1051.000000 317.850000 1056.000000 318.150000 ;
        RECT 1051.000000 325.850000 1056.000000 326.150000 ;
        RECT 1051.000000 329.850000 1056.000000 330.150000 ;
        RECT 1051.000000 333.850000 1056.000000 334.150000 ;
        RECT 1051.000000 337.850000 1056.000000 338.150000 ;
        RECT 1051.000000 341.850000 1056.000000 342.150000 ;
        RECT 1101.000000 313.850000 1106.000000 314.150000 ;
        RECT 1101.000000 309.850000 1106.000000 310.150000 ;
        RECT 1101.000000 317.850000 1106.000000 318.150000 ;
        RECT 1101.000000 321.850000 1106.000000 322.150000 ;
        RECT 1101.000000 325.850000 1106.000000 326.150000 ;
        RECT 1101.000000 329.850000 1106.000000 330.150000 ;
        RECT 1101.000000 333.850000 1106.000000 334.150000 ;
        RECT 1101.000000 337.850000 1106.000000 338.150000 ;
        RECT 1101.000000 341.850000 1106.000000 342.150000 ;
        RECT 1151.000000 305.850000 1156.000000 306.150000 ;
        RECT 1172.000000 305.850000 1182.000000 306.150000 ;
        RECT 1151.000000 277.850000 1156.000000 278.150000 ;
        RECT 1151.000000 269.850000 1156.000000 270.150000 ;
        RECT 1151.000000 273.850000 1156.000000 274.150000 ;
        RECT 1151.000000 281.850000 1156.000000 282.150000 ;
        RECT 1151.000000 285.850000 1156.000000 286.150000 ;
        RECT 1172.000000 277.850000 1182.000000 278.150000 ;
        RECT 1172.000000 269.850000 1182.000000 270.150000 ;
        RECT 1172.000000 273.850000 1182.000000 274.150000 ;
        RECT 1172.000000 281.850000 1182.000000 282.150000 ;
        RECT 1172.000000 285.850000 1182.000000 286.150000 ;
        RECT 1151.000000 301.850000 1156.000000 302.150000 ;
        RECT 1151.000000 297.850000 1156.000000 298.150000 ;
        RECT 1151.000000 289.850000 1156.000000 290.150000 ;
        RECT 1151.000000 293.850000 1156.000000 294.150000 ;
        RECT 1172.000000 301.850000 1182.000000 302.150000 ;
        RECT 1172.000000 289.850000 1182.000000 290.150000 ;
        RECT 1172.000000 293.850000 1182.000000 294.150000 ;
        RECT 1172.000000 297.850000 1182.000000 298.150000 ;
        RECT 1151.000000 321.850000 1156.000000 322.150000 ;
        RECT 1151.000000 317.850000 1156.000000 318.150000 ;
        RECT 1151.000000 309.850000 1156.000000 310.150000 ;
        RECT 1151.000000 313.850000 1156.000000 314.150000 ;
        RECT 1172.000000 321.850000 1182.000000 322.150000 ;
        RECT 1172.000000 309.850000 1182.000000 310.150000 ;
        RECT 1172.000000 313.850000 1182.000000 314.150000 ;
        RECT 1172.000000 317.850000 1182.000000 318.150000 ;
        RECT 1151.000000 329.850000 1156.000000 330.150000 ;
        RECT 1151.000000 325.850000 1156.000000 326.150000 ;
        RECT 1151.000000 333.850000 1156.000000 334.150000 ;
        RECT 1151.000000 337.850000 1156.000000 338.150000 ;
        RECT 1151.000000 341.850000 1156.000000 342.150000 ;
        RECT 1172.000000 329.850000 1182.000000 330.150000 ;
        RECT 1172.000000 325.850000 1182.000000 326.150000 ;
        RECT 1172.000000 333.850000 1182.000000 334.150000 ;
        RECT 1172.000000 337.850000 1182.000000 338.150000 ;
        RECT 1172.000000 341.850000 1182.000000 342.150000 ;
        RECT 4.000000 357.850000 14.000000 358.150000 ;
        RECT 4.000000 353.850000 14.000000 354.150000 ;
        RECT 4.000000 345.850000 14.000000 346.150000 ;
        RECT 4.000000 349.850000 14.000000 350.150000 ;
        RECT 4.000000 369.850000 14.000000 370.150000 ;
        RECT 4.000000 365.850000 14.000000 366.150000 ;
        RECT 4.000000 361.850000 14.000000 362.150000 ;
        RECT 4.000000 377.850000 14.000000 378.150000 ;
        RECT 4.000000 373.850000 14.000000 374.150000 ;
        RECT 51.000000 354.445000 56.000000 354.745000 ;
        RECT 51.000000 345.850000 56.000000 346.150000 ;
        RECT 51.000000 369.850000 56.000000 370.150000 ;
        RECT 51.000000 365.850000 56.000000 366.150000 ;
        RECT 51.000000 361.850000 56.000000 362.150000 ;
        RECT 51.000000 373.850000 56.000000 374.150000 ;
        RECT 51.000000 377.850000 56.000000 378.150000 ;
        RECT 4.000000 397.850000 14.000000 398.150000 ;
        RECT 4.000000 393.850000 14.000000 394.150000 ;
        RECT 4.000000 389.850000 14.000000 390.150000 ;
        RECT 4.000000 381.850000 14.000000 382.150000 ;
        RECT 4.000000 385.850000 14.000000 386.150000 ;
        RECT 4.000000 401.850000 14.000000 402.150000 ;
        RECT 4.000000 405.850000 14.000000 406.150000 ;
        RECT 4.000000 409.850000 14.000000 410.150000 ;
        RECT 4.000000 413.850000 14.000000 414.150000 ;
        RECT 51.000000 385.850000 56.000000 386.150000 ;
        RECT 51.000000 381.850000 56.000000 382.150000 ;
        RECT 51.000000 389.850000 56.000000 390.150000 ;
        RECT 51.000000 393.850000 56.000000 394.150000 ;
        RECT 51.000000 397.850000 56.000000 398.150000 ;
        RECT 51.000000 413.850000 56.000000 414.150000 ;
        RECT 51.000000 409.850000 56.000000 410.150000 ;
        RECT 51.000000 405.850000 56.000000 406.150000 ;
        RECT 51.000000 401.850000 56.000000 402.150000 ;
        RECT 101.000000 345.850000 106.000000 346.150000 ;
        RECT 101.000000 349.850000 106.000000 350.150000 ;
        RECT 101.000000 353.850000 106.000000 354.150000 ;
        RECT 101.000000 357.850000 106.000000 358.150000 ;
        RECT 101.000000 361.850000 106.000000 362.150000 ;
        RECT 101.000000 365.850000 106.000000 366.150000 ;
        RECT 101.000000 369.850000 106.000000 370.150000 ;
        RECT 101.000000 373.850000 106.000000 374.150000 ;
        RECT 101.000000 377.850000 106.000000 378.150000 ;
        RECT 101.000000 381.850000 106.000000 382.150000 ;
        RECT 101.000000 385.850000 106.000000 386.150000 ;
        RECT 101.000000 389.850000 106.000000 390.150000 ;
        RECT 101.000000 393.850000 106.000000 394.150000 ;
        RECT 101.000000 397.850000 106.000000 398.150000 ;
        RECT 101.000000 413.850000 106.000000 414.150000 ;
        RECT 101.000000 409.850000 106.000000 410.150000 ;
        RECT 101.000000 405.850000 106.000000 406.150000 ;
        RECT 101.000000 401.850000 106.000000 402.150000 ;
        RECT 4.000000 433.850000 14.000000 434.150000 ;
        RECT 4.000000 429.850000 14.000000 430.150000 ;
        RECT 4.000000 417.850000 14.000000 418.150000 ;
        RECT 4.000000 421.850000 14.000000 422.150000 ;
        RECT 4.000000 425.850000 14.000000 426.150000 ;
        RECT 4.000000 437.850000 14.000000 438.150000 ;
        RECT 4.000000 441.850000 14.000000 442.150000 ;
        RECT 4.000000 445.850000 14.000000 446.150000 ;
        RECT 4.000000 449.850000 14.000000 450.150000 ;
        RECT 4.000000 453.850000 14.000000 454.150000 ;
        RECT 51.000000 417.850000 56.000000 418.150000 ;
        RECT 51.000000 421.850000 56.000000 422.150000 ;
        RECT 51.000000 425.850000 56.000000 426.150000 ;
        RECT 51.000000 429.850000 56.000000 430.150000 ;
        RECT 51.000000 433.850000 56.000000 434.150000 ;
        RECT 51.000000 453.850000 56.000000 454.150000 ;
        RECT 51.000000 449.850000 56.000000 450.150000 ;
        RECT 51.000000 445.850000 56.000000 446.150000 ;
        RECT 51.000000 441.850000 56.000000 442.150000 ;
        RECT 51.000000 437.850000 56.000000 438.150000 ;
        RECT 4.000000 469.850000 14.000000 470.150000 ;
        RECT 4.000000 457.850000 14.000000 458.150000 ;
        RECT 4.000000 461.850000 14.000000 462.150000 ;
        RECT 4.000000 465.850000 14.000000 466.150000 ;
        RECT 4.000000 473.850000 14.000000 474.150000 ;
        RECT 4.000000 477.850000 14.000000 478.150000 ;
        RECT 4.000000 481.850000 14.000000 482.150000 ;
        RECT 4.000000 485.850000 14.000000 486.150000 ;
        RECT 4.000000 489.850000 14.000000 490.150000 ;
        RECT 51.000000 461.850000 56.000000 462.150000 ;
        RECT 51.000000 457.850000 56.000000 458.150000 ;
        RECT 51.000000 465.850000 56.000000 466.150000 ;
        RECT 51.000000 469.850000 56.000000 470.150000 ;
        RECT 51.000000 489.850000 56.000000 490.150000 ;
        RECT 51.000000 485.850000 56.000000 486.150000 ;
        RECT 51.000000 481.850000 56.000000 482.150000 ;
        RECT 51.000000 477.850000 56.000000 478.150000 ;
        RECT 51.000000 473.850000 56.000000 474.150000 ;
        RECT 101.000000 417.850000 106.000000 418.150000 ;
        RECT 101.000000 421.850000 106.000000 422.150000 ;
        RECT 101.000000 425.850000 106.000000 426.150000 ;
        RECT 101.000000 429.850000 106.000000 430.150000 ;
        RECT 101.000000 433.850000 106.000000 434.150000 ;
        RECT 101.000000 437.850000 106.000000 438.150000 ;
        RECT 101.000000 441.850000 106.000000 442.150000 ;
        RECT 101.000000 445.850000 106.000000 446.150000 ;
        RECT 101.000000 449.850000 106.000000 450.150000 ;
        RECT 101.000000 453.850000 106.000000 454.150000 ;
        RECT 101.000000 469.850000 106.000000 470.150000 ;
        RECT 101.000000 465.850000 106.000000 466.150000 ;
        RECT 101.000000 461.850000 106.000000 462.150000 ;
        RECT 101.000000 457.850000 106.000000 458.150000 ;
        RECT 101.000000 473.850000 106.000000 474.150000 ;
        RECT 101.000000 477.850000 106.000000 478.150000 ;
        RECT 101.000000 481.850000 106.000000 482.150000 ;
        RECT 101.000000 485.850000 106.000000 486.150000 ;
        RECT 101.000000 489.850000 106.000000 490.150000 ;
        RECT 151.000000 349.850000 156.000000 350.150000 ;
        RECT 151.000000 345.850000 156.000000 346.150000 ;
        RECT 151.000000 353.850000 156.000000 354.150000 ;
        RECT 151.000000 357.850000 156.000000 358.150000 ;
        RECT 151.000000 361.850000 156.000000 362.150000 ;
        RECT 151.000000 365.850000 156.000000 366.150000 ;
        RECT 151.000000 369.850000 156.000000 370.150000 ;
        RECT 151.000000 373.850000 156.000000 374.150000 ;
        RECT 151.000000 377.850000 156.000000 378.150000 ;
        RECT 201.000000 349.850000 206.000000 350.150000 ;
        RECT 201.000000 345.850000 206.000000 346.150000 ;
        RECT 201.000000 353.850000 206.000000 354.150000 ;
        RECT 201.000000 357.850000 206.000000 358.150000 ;
        RECT 201.000000 377.850000 206.000000 378.150000 ;
        RECT 201.000000 373.850000 206.000000 374.150000 ;
        RECT 201.000000 369.850000 206.000000 370.150000 ;
        RECT 201.000000 365.850000 206.000000 366.150000 ;
        RECT 201.000000 361.850000 206.000000 362.150000 ;
        RECT 151.000000 385.850000 156.000000 386.150000 ;
        RECT 151.000000 381.850000 156.000000 382.150000 ;
        RECT 151.000000 393.850000 156.000000 394.150000 ;
        RECT 151.000000 389.850000 156.000000 390.150000 ;
        RECT 151.000000 397.850000 156.000000 398.150000 ;
        RECT 151.000000 401.850000 156.000000 402.150000 ;
        RECT 201.000000 381.850000 206.000000 382.150000 ;
        RECT 201.000000 385.850000 206.000000 386.150000 ;
        RECT 201.000000 397.850000 206.000000 398.150000 ;
        RECT 201.000000 393.850000 206.000000 394.150000 ;
        RECT 201.000000 389.850000 206.000000 390.150000 ;
        RECT 201.000000 413.850000 206.000000 414.150000 ;
        RECT 201.000000 409.850000 206.000000 410.150000 ;
        RECT 201.000000 405.850000 206.000000 406.150000 ;
        RECT 201.000000 401.850000 206.000000 402.150000 ;
        RECT 251.000000 345.850000 256.000000 346.150000 ;
        RECT 251.000000 349.850000 256.000000 350.150000 ;
        RECT 251.000000 353.850000 256.000000 354.150000 ;
        RECT 251.000000 357.850000 256.000000 358.150000 ;
        RECT 251.000000 365.850000 256.000000 366.150000 ;
        RECT 251.000000 361.850000 256.000000 362.150000 ;
        RECT 251.000000 369.850000 256.000000 370.150000 ;
        RECT 251.000000 373.850000 256.000000 374.150000 ;
        RECT 251.000000 377.850000 256.000000 378.150000 ;
        RECT 251.000000 381.850000 256.000000 382.150000 ;
        RECT 251.000000 385.850000 256.000000 386.150000 ;
        RECT 251.000000 393.850000 256.000000 394.150000 ;
        RECT 251.000000 389.850000 256.000000 390.150000 ;
        RECT 251.000000 397.850000 256.000000 398.150000 ;
        RECT 251.000000 401.850000 256.000000 402.150000 ;
        RECT 151.000000 453.850000 156.000000 454.150000 ;
        RECT 201.000000 425.850000 206.000000 426.150000 ;
        RECT 201.000000 421.850000 206.000000 422.150000 ;
        RECT 201.000000 417.850000 206.000000 418.150000 ;
        RECT 201.000000 429.850000 206.000000 430.150000 ;
        RECT 201.000000 433.850000 206.000000 434.150000 ;
        RECT 201.000000 453.850000 206.000000 454.150000 ;
        RECT 201.000000 449.850000 206.000000 450.150000 ;
        RECT 201.000000 445.850000 206.000000 446.150000 ;
        RECT 201.000000 441.850000 206.000000 442.150000 ;
        RECT 201.000000 437.850000 206.000000 438.150000 ;
        RECT 151.000000 461.850000 156.000000 462.150000 ;
        RECT 151.000000 457.850000 156.000000 458.150000 ;
        RECT 151.000000 469.850000 156.000000 470.150000 ;
        RECT 151.000000 465.850000 156.000000 466.150000 ;
        RECT 151.000000 481.850000 156.000000 482.150000 ;
        RECT 151.000000 477.850000 156.000000 478.150000 ;
        RECT 151.000000 473.850000 156.000000 474.150000 ;
        RECT 151.000000 489.850000 156.000000 490.150000 ;
        RECT 151.000000 485.850000 156.000000 486.150000 ;
        RECT 201.000000 461.850000 206.000000 462.150000 ;
        RECT 201.000000 457.850000 206.000000 458.150000 ;
        RECT 201.000000 465.850000 206.000000 466.150000 ;
        RECT 201.000000 469.850000 206.000000 470.150000 ;
        RECT 201.000000 489.850000 206.000000 490.150000 ;
        RECT 201.000000 485.850000 206.000000 486.150000 ;
        RECT 201.000000 481.850000 206.000000 482.150000 ;
        RECT 201.000000 477.850000 206.000000 478.150000 ;
        RECT 201.000000 473.850000 206.000000 474.150000 ;
        RECT 251.000000 453.850000 256.000000 454.150000 ;
        RECT 251.000000 457.850000 256.000000 458.150000 ;
        RECT 251.000000 461.850000 256.000000 462.150000 ;
        RECT 251.000000 465.850000 256.000000 466.150000 ;
        RECT 251.000000 469.850000 256.000000 470.150000 ;
        RECT 251.000000 481.850000 256.000000 482.150000 ;
        RECT 251.000000 473.850000 256.000000 474.150000 ;
        RECT 251.000000 477.850000 256.000000 478.150000 ;
        RECT 251.000000 485.850000 256.000000 486.150000 ;
        RECT 251.000000 489.850000 256.000000 490.150000 ;
        RECT 4.000000 505.850000 14.000000 506.150000 ;
        RECT 4.000000 497.850000 14.000000 498.150000 ;
        RECT 4.000000 493.850000 14.000000 494.150000 ;
        RECT 4.000000 501.850000 14.000000 502.150000 ;
        RECT 4.000000 513.850000 14.000000 514.150000 ;
        RECT 4.000000 509.850000 14.000000 510.150000 ;
        RECT 51.000000 493.850000 56.000000 494.150000 ;
        RECT 51.000000 497.850000 56.000000 498.150000 ;
        RECT 51.000000 501.850000 56.000000 502.150000 ;
        RECT 51.000000 505.850000 56.000000 506.150000 ;
        RECT 51.000000 513.850000 56.000000 514.150000 ;
        RECT 51.000000 509.850000 56.000000 510.150000 ;
        RECT 101.000000 505.850000 106.000000 506.150000 ;
        RECT 101.000000 501.850000 106.000000 502.150000 ;
        RECT 101.000000 497.850000 106.000000 498.150000 ;
        RECT 101.000000 493.850000 106.000000 494.150000 ;
        RECT 101.000000 513.850000 106.000000 514.150000 ;
        RECT 101.000000 509.850000 106.000000 510.150000 ;
        RECT 151.000000 493.850000 156.000000 494.150000 ;
        RECT 151.000000 497.850000 156.000000 498.150000 ;
        RECT 151.000000 501.850000 156.000000 502.150000 ;
        RECT 151.000000 505.850000 156.000000 506.150000 ;
        RECT 151.000000 513.850000 156.000000 514.150000 ;
        RECT 151.000000 509.850000 156.000000 510.150000 ;
        RECT 201.000000 497.850000 206.000000 498.150000 ;
        RECT 201.000000 493.850000 206.000000 494.150000 ;
        RECT 201.000000 501.850000 206.000000 502.150000 ;
        RECT 201.000000 505.850000 206.000000 506.150000 ;
        RECT 201.000000 513.850000 206.000000 514.150000 ;
        RECT 201.000000 509.850000 206.000000 510.150000 ;
        RECT 251.000000 493.850000 256.000000 494.150000 ;
        RECT 251.000000 497.850000 256.000000 498.150000 ;
        RECT 251.000000 501.850000 256.000000 502.150000 ;
        RECT 251.000000 505.850000 256.000000 506.150000 ;
        RECT 251.000000 513.850000 256.000000 514.150000 ;
        RECT 251.000000 509.850000 256.000000 510.150000 ;
        RECT 301.000000 345.850000 306.000000 346.150000 ;
        RECT 301.000000 349.850000 306.000000 350.150000 ;
        RECT 301.000000 353.850000 306.000000 354.150000 ;
        RECT 301.000000 357.850000 306.000000 358.150000 ;
        RECT 301.000000 369.850000 306.000000 370.150000 ;
        RECT 301.000000 365.850000 306.000000 366.150000 ;
        RECT 301.000000 361.850000 306.000000 362.150000 ;
        RECT 301.000000 377.850000 306.000000 378.150000 ;
        RECT 301.000000 373.850000 306.000000 374.150000 ;
        RECT 351.000000 345.850000 356.000000 346.150000 ;
        RECT 351.000000 349.850000 356.000000 350.150000 ;
        RECT 351.000000 353.850000 356.000000 354.150000 ;
        RECT 351.000000 357.850000 356.000000 358.150000 ;
        RECT 351.000000 377.850000 356.000000 378.150000 ;
        RECT 351.000000 373.850000 356.000000 374.150000 ;
        RECT 351.000000 369.850000 356.000000 370.150000 ;
        RECT 351.000000 365.850000 356.000000 366.150000 ;
        RECT 351.000000 361.850000 356.000000 362.150000 ;
        RECT 301.000000 385.850000 306.000000 386.150000 ;
        RECT 301.000000 381.850000 306.000000 382.150000 ;
        RECT 301.000000 389.850000 306.000000 390.150000 ;
        RECT 301.000000 393.850000 306.000000 394.150000 ;
        RECT 301.000000 397.850000 306.000000 398.150000 ;
        RECT 301.000000 405.850000 306.000000 406.150000 ;
        RECT 301.000000 401.850000 306.000000 402.150000 ;
        RECT 301.000000 413.850000 306.000000 414.150000 ;
        RECT 301.000000 409.850000 306.000000 410.150000 ;
        RECT 351.000000 381.850000 356.000000 382.150000 ;
        RECT 351.000000 385.850000 356.000000 386.150000 ;
        RECT 351.000000 397.850000 356.000000 398.150000 ;
        RECT 351.000000 393.850000 356.000000 394.150000 ;
        RECT 351.000000 389.850000 356.000000 390.150000 ;
        RECT 351.000000 413.850000 356.000000 414.150000 ;
        RECT 351.000000 409.850000 356.000000 410.150000 ;
        RECT 351.000000 405.850000 356.000000 406.150000 ;
        RECT 351.000000 401.850000 356.000000 402.150000 ;
        RECT 401.000000 357.850000 406.000000 358.150000 ;
        RECT 401.000000 353.850000 406.000000 354.150000 ;
        RECT 401.000000 349.850000 406.000000 350.150000 ;
        RECT 401.000000 345.850000 406.000000 346.150000 ;
        RECT 401.000000 361.850000 406.000000 362.150000 ;
        RECT 401.000000 365.850000 406.000000 366.150000 ;
        RECT 401.000000 369.850000 406.000000 370.150000 ;
        RECT 401.000000 377.850000 406.000000 378.150000 ;
        RECT 401.000000 373.850000 406.000000 374.150000 ;
        RECT 401.000000 385.850000 406.000000 386.150000 ;
        RECT 401.000000 381.850000 406.000000 382.150000 ;
        RECT 401.000000 397.850000 406.000000 398.150000 ;
        RECT 401.000000 393.850000 406.000000 394.150000 ;
        RECT 401.000000 389.850000 406.000000 390.150000 ;
        RECT 401.000000 401.850000 406.000000 402.150000 ;
        RECT 401.000000 405.850000 406.000000 406.150000 ;
        RECT 401.000000 409.850000 406.000000 410.150000 ;
        RECT 401.000000 413.850000 406.000000 414.150000 ;
        RECT 301.000000 425.850000 306.000000 426.150000 ;
        RECT 301.000000 417.850000 306.000000 418.150000 ;
        RECT 301.000000 421.850000 306.000000 422.150000 ;
        RECT 301.000000 429.850000 306.000000 430.150000 ;
        RECT 301.000000 433.850000 306.000000 434.150000 ;
        RECT 301.000000 441.850000 306.000000 442.150000 ;
        RECT 301.000000 437.850000 306.000000 438.150000 ;
        RECT 301.000000 453.850000 306.000000 454.150000 ;
        RECT 301.000000 449.850000 306.000000 450.150000 ;
        RECT 301.000000 445.850000 306.000000 446.150000 ;
        RECT 351.000000 417.850000 356.000000 418.150000 ;
        RECT 351.000000 421.850000 356.000000 422.150000 ;
        RECT 351.000000 425.850000 356.000000 426.150000 ;
        RECT 351.000000 429.850000 356.000000 430.150000 ;
        RECT 351.000000 433.850000 356.000000 434.150000 ;
        RECT 351.000000 437.850000 356.000000 438.150000 ;
        RECT 351.000000 441.850000 356.000000 442.150000 ;
        RECT 351.000000 445.850000 356.000000 446.150000 ;
        RECT 351.000000 449.850000 356.000000 450.150000 ;
        RECT 351.000000 453.850000 356.000000 454.150000 ;
        RECT 301.000000 461.850000 306.000000 462.150000 ;
        RECT 301.000000 457.850000 306.000000 458.150000 ;
        RECT 301.000000 465.850000 306.000000 466.150000 ;
        RECT 301.000000 469.850000 306.000000 470.150000 ;
        RECT 301.000000 481.850000 306.000000 482.150000 ;
        RECT 301.000000 477.850000 306.000000 478.150000 ;
        RECT 301.000000 473.850000 306.000000 474.150000 ;
        RECT 301.000000 489.850000 306.000000 490.150000 ;
        RECT 301.000000 485.850000 306.000000 486.150000 ;
        RECT 351.000000 461.850000 356.000000 462.150000 ;
        RECT 351.000000 457.850000 356.000000 458.150000 ;
        RECT 351.000000 465.850000 356.000000 466.150000 ;
        RECT 351.000000 469.850000 356.000000 470.150000 ;
        RECT 351.000000 481.850000 356.000000 482.150000 ;
        RECT 351.000000 473.850000 356.000000 474.150000 ;
        RECT 351.000000 477.850000 356.000000 478.150000 ;
        RECT 351.000000 485.850000 356.000000 486.150000 ;
        RECT 351.000000 489.850000 356.000000 490.150000 ;
        RECT 401.000000 417.850000 406.000000 418.150000 ;
        RECT 401.000000 421.850000 406.000000 422.150000 ;
        RECT 401.000000 425.850000 406.000000 426.150000 ;
        RECT 401.000000 433.850000 406.000000 434.150000 ;
        RECT 401.000000 429.850000 406.000000 430.150000 ;
        RECT 401.000000 437.850000 406.000000 438.150000 ;
        RECT 401.000000 441.850000 406.000000 442.150000 ;
        RECT 401.000000 445.850000 406.000000 446.150000 ;
        RECT 401.000000 449.850000 406.000000 450.150000 ;
        RECT 401.000000 453.850000 406.000000 454.150000 ;
        RECT 401.000000 461.850000 406.000000 462.150000 ;
        RECT 401.000000 457.850000 406.000000 458.150000 ;
        RECT 401.000000 465.850000 406.000000 466.150000 ;
        RECT 401.000000 469.850000 406.000000 470.150000 ;
        RECT 401.000000 481.850000 406.000000 482.150000 ;
        RECT 401.000000 473.850000 406.000000 474.150000 ;
        RECT 401.000000 477.850000 406.000000 478.150000 ;
        RECT 401.000000 485.850000 406.000000 486.150000 ;
        RECT 401.000000 489.850000 406.000000 490.150000 ;
        RECT 451.000000 345.850000 456.000000 346.150000 ;
        RECT 451.000000 369.850000 456.000000 370.150000 ;
        RECT 451.000000 377.850000 456.000000 378.150000 ;
        RECT 451.000000 373.850000 456.000000 374.150000 ;
        RECT 451.000000 366.105000 456.000000 367.105000 ;
        RECT 501.000000 345.850000 506.000000 346.150000 ;
        RECT 501.000000 349.850000 506.000000 350.150000 ;
        RECT 501.000000 353.850000 506.000000 354.150000 ;
        RECT 501.000000 357.850000 506.000000 358.150000 ;
        RECT 501.000000 361.850000 506.000000 362.150000 ;
        RECT 501.000000 365.850000 506.000000 366.150000 ;
        RECT 501.000000 369.850000 506.000000 370.150000 ;
        RECT 501.000000 377.850000 506.000000 378.150000 ;
        RECT 501.000000 373.850000 506.000000 374.150000 ;
        RECT 451.000000 381.850000 456.000000 382.150000 ;
        RECT 451.000000 385.850000 456.000000 386.150000 ;
        RECT 451.000000 397.850000 456.000000 398.150000 ;
        RECT 451.000000 393.850000 456.000000 394.150000 ;
        RECT 451.000000 389.850000 456.000000 390.150000 ;
        RECT 451.000000 416.105000 456.000000 417.105000 ;
        RECT 501.000000 381.850000 506.000000 382.150000 ;
        RECT 501.000000 385.850000 506.000000 386.150000 ;
        RECT 501.000000 393.850000 506.000000 394.150000 ;
        RECT 501.000000 389.850000 506.000000 390.150000 ;
        RECT 501.000000 397.850000 506.000000 398.150000 ;
        RECT 501.000000 401.850000 506.000000 402.150000 ;
        RECT 501.000000 405.850000 506.000000 406.150000 ;
        RECT 501.000000 409.850000 506.000000 410.150000 ;
        RECT 501.000000 413.850000 506.000000 414.150000 ;
        RECT 551.000000 357.850000 556.000000 358.150000 ;
        RECT 551.000000 353.850000 556.000000 354.150000 ;
        RECT 551.000000 349.850000 556.000000 350.150000 ;
        RECT 551.000000 345.850000 556.000000 346.150000 ;
        RECT 551.000000 361.850000 556.000000 362.150000 ;
        RECT 551.000000 365.850000 556.000000 366.150000 ;
        RECT 551.000000 369.850000 556.000000 370.150000 ;
        RECT 551.000000 373.850000 556.000000 374.150000 ;
        RECT 551.000000 377.850000 556.000000 378.150000 ;
        RECT 551.000000 385.850000 556.000000 386.150000 ;
        RECT 551.000000 381.850000 556.000000 382.150000 ;
        RECT 551.000000 397.850000 556.000000 398.150000 ;
        RECT 551.000000 393.850000 556.000000 394.150000 ;
        RECT 551.000000 389.850000 556.000000 390.150000 ;
        RECT 551.000000 413.850000 556.000000 414.150000 ;
        RECT 551.000000 409.850000 556.000000 410.150000 ;
        RECT 551.000000 405.850000 556.000000 406.150000 ;
        RECT 551.000000 401.850000 556.000000 402.150000 ;
        RECT 451.000000 425.850000 456.000000 426.150000 ;
        RECT 451.000000 421.850000 456.000000 422.150000 ;
        RECT 451.000000 429.850000 456.000000 430.150000 ;
        RECT 451.000000 433.850000 456.000000 434.150000 ;
        RECT 451.000000 441.850000 456.000000 442.150000 ;
        RECT 451.000000 437.850000 456.000000 438.150000 ;
        RECT 451.000000 453.850000 456.000000 454.150000 ;
        RECT 451.000000 449.850000 456.000000 450.150000 ;
        RECT 451.000000 445.850000 456.000000 446.150000 ;
        RECT 501.000000 425.850000 506.000000 426.150000 ;
        RECT 501.000000 421.850000 506.000000 422.150000 ;
        RECT 501.000000 417.850000 506.000000 418.150000 ;
        RECT 501.000000 433.850000 506.000000 434.150000 ;
        RECT 501.000000 429.850000 506.000000 430.150000 ;
        RECT 501.000000 437.850000 506.000000 438.150000 ;
        RECT 501.000000 441.850000 506.000000 442.150000 ;
        RECT 501.000000 445.850000 506.000000 446.150000 ;
        RECT 501.000000 453.850000 506.000000 454.150000 ;
        RECT 501.000000 449.850000 506.000000 450.150000 ;
        RECT 451.000000 461.850000 456.000000 462.150000 ;
        RECT 451.000000 457.850000 456.000000 458.150000 ;
        RECT 451.000000 465.850000 456.000000 466.150000 ;
        RECT 451.000000 469.850000 456.000000 470.150000 ;
        RECT 451.000000 481.850000 456.000000 482.150000 ;
        RECT 451.000000 477.850000 456.000000 478.150000 ;
        RECT 451.000000 473.850000 456.000000 474.150000 ;
        RECT 451.000000 489.850000 456.000000 490.150000 ;
        RECT 451.000000 485.850000 456.000000 486.150000 ;
        RECT 501.000000 457.850000 506.000000 458.150000 ;
        RECT 501.000000 461.850000 506.000000 462.150000 ;
        RECT 501.000000 469.850000 506.000000 470.150000 ;
        RECT 501.000000 465.850000 506.000000 466.150000 ;
        RECT 501.000000 481.850000 506.000000 482.150000 ;
        RECT 501.000000 473.850000 506.000000 474.150000 ;
        RECT 501.000000 477.850000 506.000000 478.150000 ;
        RECT 501.000000 485.850000 506.000000 486.150000 ;
        RECT 501.000000 489.850000 506.000000 490.150000 ;
        RECT 551.000000 421.850000 556.000000 422.150000 ;
        RECT 551.000000 417.850000 556.000000 418.150000 ;
        RECT 551.000000 425.850000 556.000000 426.150000 ;
        RECT 551.000000 433.850000 556.000000 434.150000 ;
        RECT 551.000000 429.850000 556.000000 430.150000 ;
        RECT 551.000000 437.850000 556.000000 438.150000 ;
        RECT 551.000000 441.850000 556.000000 442.150000 ;
        RECT 551.000000 445.850000 556.000000 446.150000 ;
        RECT 551.000000 449.850000 556.000000 450.150000 ;
        RECT 551.000000 453.850000 556.000000 454.150000 ;
        RECT 551.000000 457.850000 556.000000 458.150000 ;
        RECT 551.000000 461.850000 556.000000 462.150000 ;
        RECT 551.000000 465.850000 556.000000 466.150000 ;
        RECT 551.000000 469.850000 556.000000 470.150000 ;
        RECT 551.000000 481.850000 556.000000 482.150000 ;
        RECT 551.000000 473.850000 556.000000 474.150000 ;
        RECT 551.000000 477.850000 556.000000 478.150000 ;
        RECT 551.000000 485.850000 556.000000 486.150000 ;
        RECT 551.000000 489.850000 556.000000 490.150000 ;
        RECT 301.000000 497.850000 306.000000 498.150000 ;
        RECT 301.000000 493.850000 306.000000 494.150000 ;
        RECT 301.000000 501.850000 306.000000 502.150000 ;
        RECT 301.000000 505.850000 306.000000 506.150000 ;
        RECT 301.000000 517.850000 306.000000 518.150000 ;
        RECT 301.000000 513.850000 306.000000 514.150000 ;
        RECT 301.000000 509.850000 306.000000 510.150000 ;
        RECT 351.000000 497.850000 356.000000 498.150000 ;
        RECT 351.000000 493.850000 356.000000 494.150000 ;
        RECT 351.000000 501.850000 356.000000 502.150000 ;
        RECT 351.000000 505.850000 356.000000 506.150000 ;
        RECT 351.000000 509.850000 356.000000 510.150000 ;
        RECT 351.000000 513.850000 356.000000 514.150000 ;
        RECT 351.000000 517.850000 356.000000 518.150000 ;
        RECT 351.000000 521.850000 356.000000 522.150000 ;
        RECT 351.000000 525.850000 356.000000 526.150000 ;
        RECT 351.000000 529.850000 356.000000 530.150000 ;
        RECT 351.000000 533.850000 356.000000 534.150000 ;
        RECT 351.000000 545.850000 356.000000 546.150000 ;
        RECT 351.000000 541.850000 356.000000 542.150000 ;
        RECT 351.000000 537.850000 356.000000 538.150000 ;
        RECT 351.000000 561.850000 356.000000 562.150000 ;
        RECT 351.000000 557.850000 356.000000 558.150000 ;
        RECT 351.000000 553.850000 356.000000 554.150000 ;
        RECT 351.000000 549.850000 356.000000 550.150000 ;
        RECT 385.000000 505.850000 395.000000 506.150000 ;
        RECT 385.000000 501.850000 395.000000 502.150000 ;
        RECT 385.000000 493.850000 395.000000 494.150000 ;
        RECT 385.000000 497.850000 395.000000 498.150000 ;
        RECT 401.000000 497.850000 406.000000 498.150000 ;
        RECT 401.000000 493.850000 406.000000 494.150000 ;
        RECT 401.000000 501.850000 406.000000 502.150000 ;
        RECT 385.000000 509.850000 395.000000 510.150000 ;
        RECT 385.000000 513.850000 395.000000 514.150000 ;
        RECT 385.000000 517.850000 395.000000 518.150000 ;
        RECT 385.000000 521.850000 395.000000 522.150000 ;
        RECT 385.000000 525.850000 395.000000 526.150000 ;
        RECT 385.000000 545.850000 395.000000 546.150000 ;
        RECT 385.000000 541.850000 395.000000 542.150000 ;
        RECT 385.000000 537.850000 395.000000 538.150000 ;
        RECT 385.000000 533.850000 395.000000 534.150000 ;
        RECT 385.000000 529.850000 395.000000 530.150000 ;
        RECT 385.000000 561.850000 395.000000 562.150000 ;
        RECT 385.000000 557.850000 395.000000 558.150000 ;
        RECT 385.000000 553.850000 395.000000 554.150000 ;
        RECT 385.000000 549.850000 395.000000 550.150000 ;
        RECT 351.000000 565.850000 356.000000 566.150000 ;
        RECT 351.000000 569.850000 356.000000 570.150000 ;
        RECT 351.000000 573.850000 356.000000 574.150000 ;
        RECT 351.000000 577.850000 356.000000 578.150000 ;
        RECT 351.000000 581.850000 356.000000 582.150000 ;
        RECT 351.000000 601.850000 356.000000 602.150000 ;
        RECT 351.000000 597.850000 356.000000 598.150000 ;
        RECT 351.000000 593.850000 356.000000 594.150000 ;
        RECT 351.000000 589.850000 356.000000 590.150000 ;
        RECT 351.000000 585.850000 356.000000 586.150000 ;
        RECT 351.000000 609.850000 356.000000 610.150000 ;
        RECT 351.000000 605.850000 356.000000 606.150000 ;
        RECT 351.000000 613.850000 356.000000 614.150000 ;
        RECT 351.000000 617.850000 356.000000 618.150000 ;
        RECT 351.000000 621.850000 356.000000 622.150000 ;
        RECT 351.000000 625.850000 356.000000 626.150000 ;
        RECT 351.000000 629.850000 356.000000 630.150000 ;
        RECT 351.000000 633.850000 356.000000 634.150000 ;
        RECT 351.000000 637.850000 356.000000 638.150000 ;
        RECT 385.000000 565.850000 395.000000 566.150000 ;
        RECT 385.000000 569.850000 395.000000 570.150000 ;
        RECT 385.000000 573.850000 395.000000 574.150000 ;
        RECT 385.000000 577.850000 395.000000 578.150000 ;
        RECT 385.000000 581.850000 395.000000 582.150000 ;
        RECT 385.000000 601.850000 395.000000 602.150000 ;
        RECT 385.000000 597.850000 395.000000 598.150000 ;
        RECT 385.000000 593.850000 395.000000 594.150000 ;
        RECT 385.000000 589.850000 395.000000 590.150000 ;
        RECT 385.000000 585.850000 395.000000 586.150000 ;
        RECT 385.000000 617.850000 395.000000 618.150000 ;
        RECT 385.000000 613.850000 395.000000 614.150000 ;
        RECT 385.000000 609.850000 395.000000 610.150000 ;
        RECT 385.000000 605.850000 395.000000 606.150000 ;
        RECT 385.000000 637.850000 395.000000 638.150000 ;
        RECT 385.000000 633.850000 395.000000 634.150000 ;
        RECT 385.000000 629.850000 395.000000 630.150000 ;
        RECT 385.000000 625.850000 395.000000 626.150000 ;
        RECT 385.000000 621.850000 395.000000 622.150000 ;
        RECT 451.000000 493.850000 456.000000 494.150000 ;
        RECT 451.000000 497.850000 456.000000 498.150000 ;
        RECT 451.000000 501.850000 456.000000 502.150000 ;
        RECT 501.000000 493.850000 506.000000 494.150000 ;
        RECT 501.000000 497.850000 506.000000 498.150000 ;
        RECT 501.000000 501.850000 506.000000 502.150000 ;
        RECT 551.000000 493.850000 556.000000 494.150000 ;
        RECT 551.000000 497.850000 556.000000 498.150000 ;
        RECT 551.000000 501.850000 556.000000 502.150000 ;
        RECT 351.000000 657.850000 356.000000 658.150000 ;
        RECT 351.000000 641.850000 356.000000 642.150000 ;
        RECT 351.000000 645.850000 356.000000 646.150000 ;
        RECT 351.000000 649.850000 356.000000 650.150000 ;
        RECT 351.000000 653.850000 356.000000 654.150000 ;
        RECT 351.000000 673.850000 356.000000 674.150000 ;
        RECT 351.000000 669.850000 356.000000 670.150000 ;
        RECT 351.000000 665.850000 356.000000 666.150000 ;
        RECT 351.000000 661.850000 356.000000 662.150000 ;
        RECT 301.000000 681.850000 306.000000 682.150000 ;
        RECT 301.000000 677.850000 306.000000 678.150000 ;
        RECT 351.000000 677.850000 356.000000 678.150000 ;
        RECT 351.000000 681.850000 356.000000 682.150000 ;
        RECT 385.000000 657.850000 395.000000 658.150000 ;
        RECT 401.000000 657.850000 406.000000 658.150000 ;
        RECT 385.000000 641.850000 395.000000 642.150000 ;
        RECT 385.000000 645.850000 395.000000 646.150000 ;
        RECT 385.000000 649.850000 395.000000 650.150000 ;
        RECT 385.000000 653.850000 395.000000 654.150000 ;
        RECT 385.000000 673.850000 395.000000 674.150000 ;
        RECT 385.000000 669.850000 395.000000 670.150000 ;
        RECT 385.000000 665.850000 395.000000 666.150000 ;
        RECT 385.000000 661.850000 395.000000 662.150000 ;
        RECT 401.000000 661.850000 406.000000 662.150000 ;
        RECT 401.000000 665.850000 406.000000 666.150000 ;
        RECT 401.000000 669.850000 406.000000 670.150000 ;
        RECT 401.000000 673.850000 406.000000 674.150000 ;
        RECT 401.000000 677.850000 406.000000 678.150000 ;
        RECT 385.000000 677.850000 395.000000 678.150000 ;
        RECT 401.000000 681.850000 406.000000 682.150000 ;
        RECT 385.000000 681.850000 395.000000 682.150000 ;
        RECT 451.000000 657.850000 456.000000 658.150000 ;
        RECT 451.000000 661.850000 456.000000 662.150000 ;
        RECT 451.000000 665.850000 456.000000 666.150000 ;
        RECT 451.000000 669.850000 456.000000 670.150000 ;
        RECT 451.000000 673.850000 456.000000 674.150000 ;
        RECT 501.000000 657.850000 506.000000 658.150000 ;
        RECT 501.000000 661.850000 506.000000 662.150000 ;
        RECT 501.000000 665.850000 506.000000 666.150000 ;
        RECT 501.000000 673.850000 506.000000 674.150000 ;
        RECT 501.000000 669.850000 506.000000 670.150000 ;
        RECT 451.000000 677.850000 456.000000 678.150000 ;
        RECT 451.000000 681.850000 456.000000 682.150000 ;
        RECT 501.000000 677.850000 506.000000 678.150000 ;
        RECT 501.000000 681.850000 506.000000 682.150000 ;
        RECT 551.000000 657.850000 556.000000 658.150000 ;
        RECT 551.000000 661.850000 556.000000 662.150000 ;
        RECT 551.000000 665.850000 556.000000 666.150000 ;
        RECT 551.000000 669.850000 556.000000 670.150000 ;
        RECT 551.000000 673.850000 556.000000 674.150000 ;
        RECT 551.000000 681.850000 556.000000 682.150000 ;
        RECT 551.000000 677.850000 556.000000 678.150000 ;
        RECT 735.000000 433.850000 745.000000 434.150000 ;
        RECT 735.000000 441.850000 745.000000 442.150000 ;
        RECT 735.000000 437.850000 745.000000 438.150000 ;
        RECT 735.000000 449.850000 745.000000 450.150000 ;
        RECT 735.000000 445.850000 745.000000 446.150000 ;
        RECT 735.000000 453.850000 745.000000 454.150000 ;
        RECT 735.000000 457.850000 745.000000 458.150000 ;
        RECT 735.000000 461.850000 745.000000 462.150000 ;
        RECT 735.000000 465.850000 745.000000 466.150000 ;
        RECT 735.000000 469.850000 745.000000 470.150000 ;
        RECT 735.000000 481.850000 745.000000 482.150000 ;
        RECT 735.000000 473.850000 745.000000 474.150000 ;
        RECT 735.000000 477.850000 745.000000 478.150000 ;
        RECT 735.000000 485.850000 745.000000 486.150000 ;
        RECT 735.000000 489.850000 745.000000 490.150000 ;
        RECT 601.000000 357.850000 606.000000 358.150000 ;
        RECT 601.000000 353.850000 606.000000 354.150000 ;
        RECT 601.000000 349.850000 606.000000 350.150000 ;
        RECT 601.000000 345.850000 606.000000 346.150000 ;
        RECT 601.000000 361.850000 606.000000 362.150000 ;
        RECT 601.000000 365.850000 606.000000 366.150000 ;
        RECT 601.000000 369.850000 606.000000 370.150000 ;
        RECT 601.000000 373.850000 606.000000 374.150000 ;
        RECT 601.000000 377.850000 606.000000 378.150000 ;
        RECT 651.000000 349.850000 656.000000 350.150000 ;
        RECT 651.000000 345.850000 656.000000 346.150000 ;
        RECT 651.000000 353.850000 656.000000 354.150000 ;
        RECT 651.000000 357.850000 656.000000 358.150000 ;
        RECT 651.000000 361.850000 656.000000 362.150000 ;
        RECT 651.000000 365.850000 656.000000 366.150000 ;
        RECT 651.000000 369.850000 656.000000 370.150000 ;
        RECT 651.000000 373.850000 656.000000 374.150000 ;
        RECT 651.000000 377.850000 656.000000 378.150000 ;
        RECT 601.000000 385.850000 606.000000 386.150000 ;
        RECT 601.000000 381.850000 606.000000 382.150000 ;
        RECT 601.000000 389.850000 606.000000 390.150000 ;
        RECT 601.000000 393.850000 606.000000 394.150000 ;
        RECT 601.000000 397.850000 606.000000 398.150000 ;
        RECT 601.000000 405.850000 606.000000 406.150000 ;
        RECT 601.000000 401.850000 606.000000 402.150000 ;
        RECT 601.000000 413.850000 606.000000 414.150000 ;
        RECT 601.000000 409.850000 606.000000 410.150000 ;
        RECT 651.000000 381.850000 656.000000 382.150000 ;
        RECT 651.000000 385.850000 656.000000 386.150000 ;
        RECT 651.000000 393.850000 656.000000 394.150000 ;
        RECT 651.000000 389.850000 656.000000 390.150000 ;
        RECT 651.000000 397.850000 656.000000 398.150000 ;
        RECT 651.000000 401.850000 656.000000 402.150000 ;
        RECT 651.000000 405.850000 656.000000 406.150000 ;
        RECT 651.000000 409.850000 656.000000 410.150000 ;
        RECT 651.000000 413.850000 656.000000 414.150000 ;
        RECT 701.000000 357.850000 706.000000 358.150000 ;
        RECT 701.000000 353.850000 706.000000 354.150000 ;
        RECT 701.000000 349.850000 706.000000 350.150000 ;
        RECT 701.000000 345.850000 706.000000 346.150000 ;
        RECT 701.000000 361.850000 706.000000 362.150000 ;
        RECT 701.000000 365.850000 706.000000 366.150000 ;
        RECT 701.000000 369.850000 706.000000 370.150000 ;
        RECT 701.000000 373.850000 706.000000 374.150000 ;
        RECT 701.000000 377.850000 706.000000 378.150000 ;
        RECT 701.000000 385.850000 706.000000 386.150000 ;
        RECT 701.000000 381.850000 706.000000 382.150000 ;
        RECT 701.000000 397.850000 706.000000 398.150000 ;
        RECT 701.000000 393.850000 706.000000 394.150000 ;
        RECT 701.000000 389.850000 706.000000 390.150000 ;
        RECT 701.000000 413.850000 706.000000 414.150000 ;
        RECT 701.000000 409.850000 706.000000 410.150000 ;
        RECT 701.000000 405.850000 706.000000 406.150000 ;
        RECT 701.000000 401.850000 706.000000 402.150000 ;
        RECT 601.000000 417.850000 606.000000 418.150000 ;
        RECT 601.000000 421.850000 606.000000 422.150000 ;
        RECT 601.000000 425.850000 606.000000 426.150000 ;
        RECT 601.000000 429.850000 606.000000 430.150000 ;
        RECT 601.000000 433.850000 606.000000 434.150000 ;
        RECT 601.000000 441.850000 606.000000 442.150000 ;
        RECT 601.000000 437.850000 606.000000 438.150000 ;
        RECT 601.000000 453.850000 606.000000 454.150000 ;
        RECT 601.000000 449.850000 606.000000 450.150000 ;
        RECT 601.000000 445.850000 606.000000 446.150000 ;
        RECT 651.000000 417.850000 656.000000 418.150000 ;
        RECT 651.000000 425.850000 656.000000 426.150000 ;
        RECT 651.000000 421.850000 656.000000 422.150000 ;
        RECT 651.000000 429.850000 656.000000 430.150000 ;
        RECT 651.000000 433.850000 656.000000 434.150000 ;
        RECT 651.000000 437.850000 656.000000 438.150000 ;
        RECT 651.000000 441.850000 656.000000 442.150000 ;
        RECT 651.000000 445.850000 656.000000 446.150000 ;
        RECT 651.000000 449.850000 656.000000 450.150000 ;
        RECT 651.000000 453.850000 656.000000 454.150000 ;
        RECT 601.000000 461.850000 606.000000 462.150000 ;
        RECT 601.000000 457.850000 606.000000 458.150000 ;
        RECT 601.000000 465.850000 606.000000 466.150000 ;
        RECT 601.000000 469.850000 606.000000 470.150000 ;
        RECT 601.000000 481.850000 606.000000 482.150000 ;
        RECT 601.000000 477.850000 606.000000 478.150000 ;
        RECT 601.000000 473.850000 606.000000 474.150000 ;
        RECT 601.000000 489.850000 606.000000 490.150000 ;
        RECT 601.000000 485.850000 606.000000 486.150000 ;
        RECT 651.000000 457.850000 656.000000 458.150000 ;
        RECT 651.000000 461.850000 656.000000 462.150000 ;
        RECT 651.000000 469.850000 656.000000 470.150000 ;
        RECT 651.000000 465.850000 656.000000 466.150000 ;
        RECT 651.000000 481.850000 656.000000 482.150000 ;
        RECT 651.000000 477.850000 656.000000 478.150000 ;
        RECT 651.000000 473.850000 656.000000 474.150000 ;
        RECT 651.000000 489.850000 656.000000 490.150000 ;
        RECT 651.000000 485.850000 656.000000 486.150000 ;
        RECT 701.000000 417.850000 706.000000 418.150000 ;
        RECT 701.000000 421.850000 706.000000 422.150000 ;
        RECT 701.000000 425.850000 706.000000 426.150000 ;
        RECT 701.000000 433.850000 706.000000 434.150000 ;
        RECT 701.000000 429.850000 706.000000 430.150000 ;
        RECT 701.000000 437.850000 706.000000 438.150000 ;
        RECT 701.000000 441.850000 706.000000 442.150000 ;
        RECT 701.000000 445.850000 706.000000 446.150000 ;
        RECT 701.000000 449.850000 706.000000 450.150000 ;
        RECT 701.000000 453.850000 706.000000 454.150000 ;
        RECT 701.000000 457.850000 706.000000 458.150000 ;
        RECT 701.000000 461.850000 706.000000 462.150000 ;
        RECT 701.000000 465.850000 706.000000 466.150000 ;
        RECT 701.000000 469.850000 706.000000 470.150000 ;
        RECT 701.000000 481.850000 706.000000 482.150000 ;
        RECT 701.000000 473.850000 706.000000 474.150000 ;
        RECT 701.000000 477.850000 706.000000 478.150000 ;
        RECT 701.000000 485.850000 706.000000 486.150000 ;
        RECT 701.000000 489.850000 706.000000 490.150000 ;
        RECT 751.000000 357.850000 756.000000 358.150000 ;
        RECT 751.000000 353.850000 756.000000 354.150000 ;
        RECT 751.000000 349.850000 756.000000 350.150000 ;
        RECT 751.000000 345.850000 756.000000 346.150000 ;
        RECT 751.000000 361.850000 756.000000 362.150000 ;
        RECT 751.000000 365.850000 756.000000 366.150000 ;
        RECT 751.000000 369.850000 756.000000 370.150000 ;
        RECT 751.000000 373.850000 756.000000 374.150000 ;
        RECT 751.000000 377.850000 756.000000 378.150000 ;
        RECT 801.000000 349.850000 806.000000 350.150000 ;
        RECT 801.000000 345.850000 806.000000 346.150000 ;
        RECT 801.000000 353.850000 806.000000 354.150000 ;
        RECT 801.000000 357.850000 806.000000 358.150000 ;
        RECT 801.000000 361.850000 806.000000 362.150000 ;
        RECT 801.000000 365.850000 806.000000 366.150000 ;
        RECT 801.000000 369.850000 806.000000 370.150000 ;
        RECT 801.000000 377.850000 806.000000 378.150000 ;
        RECT 801.000000 373.850000 806.000000 374.150000 ;
        RECT 751.000000 385.850000 756.000000 386.150000 ;
        RECT 751.000000 381.850000 756.000000 382.150000 ;
        RECT 751.000000 393.850000 756.000000 394.150000 ;
        RECT 751.000000 389.850000 756.000000 390.150000 ;
        RECT 751.000000 397.850000 756.000000 398.150000 ;
        RECT 751.000000 401.850000 756.000000 402.150000 ;
        RECT 751.000000 405.850000 756.000000 406.150000 ;
        RECT 751.000000 413.850000 756.000000 414.150000 ;
        RECT 751.000000 409.850000 756.000000 410.150000 ;
        RECT 801.000000 385.850000 806.000000 386.150000 ;
        RECT 801.000000 381.850000 806.000000 382.150000 ;
        RECT 801.000000 393.850000 806.000000 394.150000 ;
        RECT 801.000000 389.850000 806.000000 390.150000 ;
        RECT 801.000000 397.850000 806.000000 398.150000 ;
        RECT 801.000000 401.850000 806.000000 402.150000 ;
        RECT 801.000000 405.850000 806.000000 406.150000 ;
        RECT 801.000000 413.850000 806.000000 414.150000 ;
        RECT 801.000000 409.850000 806.000000 410.150000 ;
        RECT 851.000000 357.850000 856.000000 358.150000 ;
        RECT 851.000000 353.850000 856.000000 354.150000 ;
        RECT 851.000000 349.850000 856.000000 350.150000 ;
        RECT 851.000000 345.850000 856.000000 346.150000 ;
        RECT 851.000000 361.850000 856.000000 362.150000 ;
        RECT 851.000000 365.850000 856.000000 366.150000 ;
        RECT 851.000000 369.850000 856.000000 370.150000 ;
        RECT 851.000000 373.850000 856.000000 374.150000 ;
        RECT 851.000000 377.850000 856.000000 378.150000 ;
        RECT 851.000000 385.850000 856.000000 386.150000 ;
        RECT 851.000000 381.850000 856.000000 382.150000 ;
        RECT 851.000000 397.850000 856.000000 398.150000 ;
        RECT 851.000000 393.850000 856.000000 394.150000 ;
        RECT 851.000000 389.850000 856.000000 390.150000 ;
        RECT 851.000000 413.850000 856.000000 414.150000 ;
        RECT 851.000000 409.850000 856.000000 410.150000 ;
        RECT 851.000000 405.850000 856.000000 406.150000 ;
        RECT 851.000000 401.850000 856.000000 402.150000 ;
        RECT 751.000000 417.850000 756.000000 418.150000 ;
        RECT 751.000000 421.850000 756.000000 422.150000 ;
        RECT 751.000000 425.850000 756.000000 426.150000 ;
        RECT 751.000000 429.850000 756.000000 430.150000 ;
        RECT 751.000000 433.850000 756.000000 434.150000 ;
        RECT 751.000000 437.850000 756.000000 438.150000 ;
        RECT 751.000000 441.850000 756.000000 442.150000 ;
        RECT 801.000000 417.850000 806.000000 418.150000 ;
        RECT 801.000000 421.850000 806.000000 422.150000 ;
        RECT 801.000000 425.850000 806.000000 426.150000 ;
        RECT 801.000000 433.850000 806.000000 434.150000 ;
        RECT 801.000000 429.850000 806.000000 430.150000 ;
        RECT 801.000000 437.850000 806.000000 438.150000 ;
        RECT 801.000000 441.850000 806.000000 442.150000 ;
        RECT 851.000000 433.850000 856.000000 434.150000 ;
        RECT 851.000000 429.850000 856.000000 430.150000 ;
        RECT 851.000000 425.850000 856.000000 426.150000 ;
        RECT 851.000000 421.850000 856.000000 422.150000 ;
        RECT 851.000000 417.850000 856.000000 418.150000 ;
        RECT 851.000000 441.850000 856.000000 442.150000 ;
        RECT 851.000000 437.850000 856.000000 438.150000 ;
        RECT 735.000000 501.850000 745.000000 502.150000 ;
        RECT 735.000000 497.850000 745.000000 498.150000 ;
        RECT 735.000000 493.850000 745.000000 494.150000 ;
        RECT 601.000000 501.850000 606.000000 502.150000 ;
        RECT 601.000000 493.850000 606.000000 494.150000 ;
        RECT 601.000000 497.850000 606.000000 498.150000 ;
        RECT 651.000000 497.850000 656.000000 498.150000 ;
        RECT 651.000000 493.850000 656.000000 494.150000 ;
        RECT 651.000000 501.850000 656.000000 502.150000 ;
        RECT 701.000000 493.850000 706.000000 494.150000 ;
        RECT 701.000000 497.850000 706.000000 498.150000 ;
        RECT 701.000000 501.850000 706.000000 502.150000 ;
        RECT 901.000000 357.850000 906.000000 358.150000 ;
        RECT 901.000000 353.850000 906.000000 354.150000 ;
        RECT 901.000000 349.850000 906.000000 350.150000 ;
        RECT 901.000000 345.850000 906.000000 346.150000 ;
        RECT 901.000000 361.850000 906.000000 362.150000 ;
        RECT 901.000000 365.850000 906.000000 366.150000 ;
        RECT 901.000000 369.850000 906.000000 370.150000 ;
        RECT 901.000000 373.850000 906.000000 374.150000 ;
        RECT 901.000000 377.850000 906.000000 378.150000 ;
        RECT 951.000000 345.850000 956.000000 346.150000 ;
        RECT 951.000000 349.850000 956.000000 350.150000 ;
        RECT 951.000000 353.850000 956.000000 354.150000 ;
        RECT 951.000000 357.850000 956.000000 358.150000 ;
        RECT 951.000000 361.850000 956.000000 362.150000 ;
        RECT 951.000000 365.850000 956.000000 366.150000 ;
        RECT 951.000000 369.850000 956.000000 370.150000 ;
        RECT 951.000000 373.850000 956.000000 374.150000 ;
        RECT 951.000000 377.850000 956.000000 378.150000 ;
        RECT 901.000000 385.850000 906.000000 386.150000 ;
        RECT 901.000000 381.850000 906.000000 382.150000 ;
        RECT 901.000000 393.850000 906.000000 394.150000 ;
        RECT 901.000000 389.850000 906.000000 390.150000 ;
        RECT 901.000000 397.850000 906.000000 398.150000 ;
        RECT 901.000000 401.850000 906.000000 402.150000 ;
        RECT 901.000000 405.850000 906.000000 406.150000 ;
        RECT 901.000000 413.850000 906.000000 414.150000 ;
        RECT 901.000000 409.850000 906.000000 410.150000 ;
        RECT 951.000000 385.850000 956.000000 386.150000 ;
        RECT 951.000000 381.850000 956.000000 382.150000 ;
        RECT 951.000000 389.850000 956.000000 390.150000 ;
        RECT 951.000000 393.850000 956.000000 394.150000 ;
        RECT 951.000000 397.850000 956.000000 398.150000 ;
        RECT 951.000000 405.850000 956.000000 406.150000 ;
        RECT 951.000000 401.850000 956.000000 402.150000 ;
        RECT 951.000000 413.850000 956.000000 414.150000 ;
        RECT 951.000000 409.850000 956.000000 410.150000 ;
        RECT 1001.000000 349.850000 1006.000000 350.150000 ;
        RECT 1001.000000 345.850000 1006.000000 346.150000 ;
        RECT 1001.000000 353.850000 1006.000000 354.150000 ;
        RECT 1001.000000 357.850000 1006.000000 358.150000 ;
        RECT 1001.000000 361.850000 1006.000000 362.150000 ;
        RECT 1001.000000 365.850000 1006.000000 366.150000 ;
        RECT 1001.000000 369.850000 1006.000000 370.150000 ;
        RECT 1001.000000 377.850000 1006.000000 378.150000 ;
        RECT 1001.000000 373.850000 1006.000000 374.150000 ;
        RECT 1001.000000 385.850000 1006.000000 386.150000 ;
        RECT 1001.000000 381.850000 1006.000000 382.150000 ;
        RECT 1001.000000 393.850000 1006.000000 394.150000 ;
        RECT 1001.000000 389.850000 1006.000000 390.150000 ;
        RECT 1001.000000 397.850000 1006.000000 398.150000 ;
        RECT 1001.000000 405.850000 1006.000000 406.150000 ;
        RECT 1001.000000 401.850000 1006.000000 402.150000 ;
        RECT 1001.000000 413.850000 1006.000000 414.150000 ;
        RECT 1001.000000 409.850000 1006.000000 410.150000 ;
        RECT 901.000000 417.850000 906.000000 418.150000 ;
        RECT 901.000000 425.850000 906.000000 426.150000 ;
        RECT 901.000000 421.850000 906.000000 422.150000 ;
        RECT 901.000000 433.850000 906.000000 434.150000 ;
        RECT 901.000000 429.850000 906.000000 430.150000 ;
        RECT 901.000000 437.850000 906.000000 438.150000 ;
        RECT 901.000000 441.850000 906.000000 442.150000 ;
        RECT 951.000000 417.850000 956.000000 418.150000 ;
        RECT 951.000000 421.850000 956.000000 422.150000 ;
        RECT 951.000000 425.850000 956.000000 426.150000 ;
        RECT 951.000000 429.850000 956.000000 430.150000 ;
        RECT 951.000000 433.850000 956.000000 434.150000 ;
        RECT 951.000000 441.850000 956.000000 442.150000 ;
        RECT 951.000000 437.850000 956.000000 438.150000 ;
        RECT 1001.000000 425.850000 1006.000000 426.150000 ;
        RECT 1001.000000 421.850000 1006.000000 422.150000 ;
        RECT 1001.000000 417.850000 1006.000000 418.150000 ;
        RECT 1001.000000 429.850000 1006.000000 430.150000 ;
        RECT 1001.000000 433.850000 1006.000000 434.150000 ;
        RECT 1001.000000 437.850000 1006.000000 438.150000 ;
        RECT 1001.000000 441.850000 1006.000000 442.150000 ;
        RECT 1051.000000 357.850000 1056.000000 358.150000 ;
        RECT 1051.000000 353.850000 1056.000000 354.150000 ;
        RECT 1051.000000 349.850000 1056.000000 350.150000 ;
        RECT 1051.000000 345.850000 1056.000000 346.150000 ;
        RECT 1051.000000 361.850000 1056.000000 362.150000 ;
        RECT 1051.000000 365.850000 1056.000000 366.150000 ;
        RECT 1051.000000 369.850000 1056.000000 370.150000 ;
        RECT 1051.000000 373.850000 1056.000000 374.150000 ;
        RECT 1051.000000 377.850000 1056.000000 378.150000 ;
        RECT 1101.000000 345.850000 1106.000000 346.150000 ;
        RECT 1101.000000 349.850000 1106.000000 350.150000 ;
        RECT 1101.000000 353.850000 1106.000000 354.150000 ;
        RECT 1101.000000 357.850000 1106.000000 358.150000 ;
        RECT 1101.000000 361.850000 1106.000000 362.150000 ;
        RECT 1101.000000 365.850000 1106.000000 366.150000 ;
        RECT 1101.000000 369.850000 1106.000000 370.150000 ;
        RECT 1101.000000 373.850000 1106.000000 374.150000 ;
        RECT 1101.000000 377.850000 1106.000000 378.150000 ;
        RECT 1051.000000 385.850000 1056.000000 386.150000 ;
        RECT 1051.000000 381.850000 1056.000000 382.150000 ;
        RECT 1051.000000 393.850000 1056.000000 394.150000 ;
        RECT 1051.000000 389.850000 1056.000000 390.150000 ;
        RECT 1051.000000 397.850000 1056.000000 398.150000 ;
        RECT 1051.000000 401.850000 1056.000000 402.150000 ;
        RECT 1051.000000 405.850000 1056.000000 406.150000 ;
        RECT 1051.000000 413.850000 1056.000000 414.150000 ;
        RECT 1051.000000 409.850000 1056.000000 410.150000 ;
        RECT 1101.000000 385.850000 1106.000000 386.150000 ;
        RECT 1101.000000 381.850000 1106.000000 382.150000 ;
        RECT 1101.000000 389.850000 1106.000000 390.150000 ;
        RECT 1101.000000 393.850000 1106.000000 394.150000 ;
        RECT 1101.000000 397.850000 1106.000000 398.150000 ;
        RECT 1101.000000 405.850000 1106.000000 406.150000 ;
        RECT 1101.000000 401.850000 1106.000000 402.150000 ;
        RECT 1101.000000 413.850000 1106.000000 414.150000 ;
        RECT 1101.000000 409.850000 1106.000000 410.150000 ;
        RECT 1151.000000 357.850000 1156.000000 358.150000 ;
        RECT 1151.000000 353.850000 1156.000000 354.150000 ;
        RECT 1151.000000 349.850000 1156.000000 350.150000 ;
        RECT 1151.000000 345.850000 1156.000000 346.150000 ;
        RECT 1172.000000 357.850000 1182.000000 358.150000 ;
        RECT 1172.000000 353.850000 1182.000000 354.150000 ;
        RECT 1172.000000 349.850000 1182.000000 350.150000 ;
        RECT 1172.000000 345.850000 1182.000000 346.150000 ;
        RECT 1151.000000 365.850000 1156.000000 366.150000 ;
        RECT 1151.000000 361.850000 1156.000000 362.150000 ;
        RECT 1151.000000 369.850000 1156.000000 370.150000 ;
        RECT 1151.000000 373.850000 1156.000000 374.150000 ;
        RECT 1151.000000 377.850000 1156.000000 378.150000 ;
        RECT 1172.000000 369.850000 1182.000000 370.150000 ;
        RECT 1172.000000 365.850000 1182.000000 366.150000 ;
        RECT 1172.000000 361.850000 1182.000000 362.150000 ;
        RECT 1172.000000 373.850000 1182.000000 374.150000 ;
        RECT 1172.000000 377.850000 1182.000000 378.150000 ;
        RECT 1151.000000 385.850000 1156.000000 386.150000 ;
        RECT 1151.000000 381.850000 1156.000000 382.150000 ;
        RECT 1151.000000 389.850000 1156.000000 390.150000 ;
        RECT 1151.000000 393.850000 1156.000000 394.150000 ;
        RECT 1151.000000 397.850000 1156.000000 398.150000 ;
        RECT 1172.000000 385.850000 1182.000000 386.150000 ;
        RECT 1172.000000 381.850000 1182.000000 382.150000 ;
        RECT 1172.000000 389.850000 1182.000000 390.150000 ;
        RECT 1172.000000 393.850000 1182.000000 394.150000 ;
        RECT 1172.000000 397.850000 1182.000000 398.150000 ;
        RECT 1151.000000 405.850000 1156.000000 406.150000 ;
        RECT 1151.000000 401.850000 1156.000000 402.150000 ;
        RECT 1151.000000 409.850000 1156.000000 410.150000 ;
        RECT 1151.000000 413.850000 1156.000000 414.150000 ;
        RECT 1172.000000 405.850000 1182.000000 406.150000 ;
        RECT 1172.000000 401.850000 1182.000000 402.150000 ;
        RECT 1172.000000 409.850000 1182.000000 410.150000 ;
        RECT 1172.000000 413.850000 1182.000000 414.150000 ;
        RECT 1051.000000 425.850000 1056.000000 426.150000 ;
        RECT 1051.000000 417.850000 1056.000000 418.150000 ;
        RECT 1051.000000 421.850000 1056.000000 422.150000 ;
        RECT 1051.000000 429.850000 1056.000000 430.150000 ;
        RECT 1051.000000 433.850000 1056.000000 434.150000 ;
        RECT 1051.000000 437.850000 1056.000000 438.150000 ;
        RECT 1051.000000 441.850000 1056.000000 442.150000 ;
        RECT 1101.000000 433.850000 1106.000000 434.150000 ;
        RECT 1101.000000 429.850000 1106.000000 430.150000 ;
        RECT 1101.000000 425.850000 1106.000000 426.150000 ;
        RECT 1101.000000 421.850000 1106.000000 422.150000 ;
        RECT 1101.000000 417.850000 1106.000000 418.150000 ;
        RECT 1101.000000 441.850000 1106.000000 442.150000 ;
        RECT 1101.000000 437.850000 1106.000000 438.150000 ;
        RECT 1151.000000 417.850000 1156.000000 418.150000 ;
        RECT 1151.000000 421.850000 1156.000000 422.150000 ;
        RECT 1151.000000 425.850000 1156.000000 426.150000 ;
        RECT 1151.000000 429.850000 1156.000000 430.150000 ;
        RECT 1151.000000 433.850000 1156.000000 434.150000 ;
        RECT 1172.000000 425.850000 1182.000000 426.150000 ;
        RECT 1172.000000 417.850000 1182.000000 418.150000 ;
        RECT 1172.000000 421.850000 1182.000000 422.150000 ;
        RECT 1172.000000 429.850000 1182.000000 430.150000 ;
        RECT 1172.000000 433.850000 1182.000000 434.150000 ;
        RECT 1151.000000 437.850000 1156.000000 438.150000 ;
        RECT 1151.000000 441.850000 1156.000000 442.150000 ;
        RECT 1151.000000 453.850000 1156.000000 454.150000 ;
        RECT 1151.000000 449.850000 1156.000000 450.150000 ;
        RECT 1151.000000 445.850000 1156.000000 446.150000 ;
        RECT 1172.000000 437.850000 1182.000000 438.150000 ;
        RECT 1172.000000 441.850000 1182.000000 442.150000 ;
        RECT 1151.000000 461.850000 1156.000000 462.150000 ;
        RECT 1151.000000 457.850000 1156.000000 458.150000 ;
        RECT 1151.000000 465.850000 1156.000000 466.150000 ;
        RECT 1151.000000 469.850000 1156.000000 470.150000 ;
        RECT 1151.000000 481.850000 1156.000000 482.150000 ;
        RECT 1151.000000 477.850000 1156.000000 478.150000 ;
        RECT 1151.000000 473.850000 1156.000000 474.150000 ;
        RECT 1151.000000 489.850000 1156.000000 490.150000 ;
        RECT 1151.000000 485.850000 1156.000000 486.150000 ;
        RECT 1151.000000 493.850000 1156.000000 494.150000 ;
        RECT 1151.000000 497.850000 1156.000000 498.150000 ;
        RECT 1151.000000 505.850000 1156.000000 506.150000 ;
        RECT 1151.000000 501.850000 1156.000000 502.150000 ;
        RECT 1151.000000 509.850000 1156.000000 510.150000 ;
        RECT 1151.000000 513.850000 1156.000000 514.150000 ;
        RECT 1151.000000 517.850000 1156.000000 518.150000 ;
        RECT 1151.000000 521.850000 1156.000000 522.150000 ;
        RECT 1151.000000 525.850000 1156.000000 526.150000 ;
        RECT 1151.000000 533.850000 1156.000000 534.150000 ;
        RECT 1151.000000 529.850000 1156.000000 530.150000 ;
        RECT 1151.000000 545.850000 1156.000000 546.150000 ;
        RECT 1151.000000 537.850000 1156.000000 538.150000 ;
        RECT 1151.000000 541.850000 1156.000000 542.150000 ;
        RECT 1151.000000 553.850000 1156.000000 554.150000 ;
        RECT 1151.000000 549.850000 1156.000000 550.150000 ;
        RECT 1151.000000 561.850000 1156.000000 562.150000 ;
        RECT 1151.000000 557.850000 1156.000000 558.150000 ;
        RECT 1151.000000 565.850000 1156.000000 566.150000 ;
        RECT 1151.000000 569.850000 1156.000000 570.150000 ;
        RECT 1151.000000 573.850000 1156.000000 574.150000 ;
        RECT 1151.000000 577.850000 1156.000000 578.150000 ;
        RECT 1151.000000 581.850000 1156.000000 582.150000 ;
        RECT 1151.000000 589.850000 1156.000000 590.150000 ;
        RECT 1151.000000 585.850000 1156.000000 586.150000 ;
        RECT 1151.000000 593.850000 1156.000000 594.150000 ;
        RECT 1151.000000 597.850000 1156.000000 598.150000 ;
        RECT 1151.000000 601.850000 1156.000000 602.150000 ;
        RECT 1151.000000 609.850000 1156.000000 610.150000 ;
        RECT 1151.000000 605.850000 1156.000000 606.150000 ;
        RECT 1151.000000 613.850000 1156.000000 614.150000 ;
        RECT 1151.000000 617.850000 1156.000000 618.150000 ;
        RECT 1151.000000 621.850000 1156.000000 622.150000 ;
        RECT 1151.000000 625.850000 1156.000000 626.150000 ;
        RECT 1151.000000 629.850000 1156.000000 630.150000 ;
        RECT 1151.000000 637.850000 1156.000000 638.150000 ;
        RECT 1151.000000 633.850000 1156.000000 634.150000 ;
        RECT 601.000000 657.850000 606.000000 658.150000 ;
        RECT 601.000000 673.850000 606.000000 674.150000 ;
        RECT 601.000000 669.850000 606.000000 670.150000 ;
        RECT 601.000000 665.850000 606.000000 666.150000 ;
        RECT 601.000000 661.850000 606.000000 662.150000 ;
        RECT 651.000000 657.850000 656.000000 658.150000 ;
        RECT 651.000000 661.850000 656.000000 662.150000 ;
        RECT 651.000000 665.850000 656.000000 666.150000 ;
        RECT 651.000000 673.850000 656.000000 674.150000 ;
        RECT 651.000000 669.850000 656.000000 670.150000 ;
        RECT 601.000000 677.850000 606.000000 678.150000 ;
        RECT 601.000000 681.850000 606.000000 682.150000 ;
        RECT 651.000000 677.850000 656.000000 678.150000 ;
        RECT 651.000000 681.850000 656.000000 682.150000 ;
        RECT 1151.000000 657.850000 1156.000000 658.150000 ;
        RECT 1151.000000 641.850000 1156.000000 642.150000 ;
        RECT 1151.000000 645.850000 1156.000000 646.150000 ;
        RECT 1151.000000 653.850000 1156.000000 654.150000 ;
        RECT 1151.000000 649.850000 1156.000000 650.150000 ;
        RECT 1151.000000 665.850000 1156.000000 666.150000 ;
        RECT 1151.000000 661.850000 1156.000000 662.150000 ;
        RECT 1151.000000 669.850000 1156.000000 670.150000 ;
        RECT 1151.000000 673.850000 1156.000000 674.150000 ;
        RECT 1151.000000 681.850000 1156.000000 682.150000 ;
        RECT 1151.000000 677.850000 1156.000000 678.150000 ;
    END
# end of P/G power stripe data as pin

  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M7 ;
        RECT 60.000000 0.000000 65.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 60.000000 681.000000 65.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 110.000000 0.000000 115.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 110.000000 681.000000 115.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 160.000000 0.000000 165.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 210.000000 0.000000 215.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 260.000000 0.000000 265.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 260.000000 681.000000 265.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 310.000000 0.000000 315.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 310.000000 681.000000 315.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 360.000000 0.000000 365.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 360.000000 681.000000 365.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 0.000000 415.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 501.000000 415.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 656.000000 415.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 410.000000 681.000000 415.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 0.000000 465.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 501.000000 465.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 656.000000 465.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 460.000000 681.000000 465.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 0.000000 515.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 501.000000 515.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 656.000000 515.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 510.000000 681.000000 515.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 0.000000 565.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 501.000000 565.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 656.000000 565.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 560.000000 681.000000 565.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 0.000000 615.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 501.000000 615.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 656.000000 615.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 610.000000 681.000000 615.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 0.000000 665.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 501.000000 665.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 656.000000 665.000000 661.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 660.000000 681.000000 665.000000 686.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 710.000000 0.000000 715.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 710.000000 501.000000 715.000000 506.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 760.000000 0.000000 765.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 760.000000 441.000000 765.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 810.000000 0.000000 815.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 810.000000 441.000000 815.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 860.000000 0.000000 865.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 860.000000 441.000000 865.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 910.000000 0.000000 915.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 910.000000 441.000000 915.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 960.000000 0.000000 965.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 960.000000 441.000000 965.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1010.000000 0.000000 1015.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1010.000000 441.000000 1015.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1060.000000 0.000000 1065.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1060.000000 441.000000 1065.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1110.000000 0.000000 1115.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1110.000000 441.000000 1115.000000 446.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1160.000000 0.000000 1165.000000 5.000000 ;
    END
    PORT
      LAYER M7 ;
        RECT 1160.000000 681.000000 1165.000000 686.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER M2 ;
        RECT 60.000000 3.850000 65.000000 4.150000 ;
        RECT 60.000000 7.850000 65.000000 8.150000 ;
        RECT 110.000000 7.850000 115.000000 8.150000 ;
        RECT 110.000000 3.850000 115.000000 4.150000 ;
        RECT 160.000000 7.850000 165.000000 8.150000 ;
        RECT 160.000000 3.850000 165.000000 4.150000 ;
        RECT 210.000000 7.850000 215.000000 8.150000 ;
        RECT 210.000000 3.850000 215.000000 4.150000 ;
        RECT 260.000000 7.850000 265.000000 8.150000 ;
        RECT 260.000000 3.850000 265.000000 4.150000 ;
        RECT 310.000000 7.850000 315.000000 8.150000 ;
        RECT 310.000000 3.850000 315.000000 4.150000 ;
        RECT 360.000000 7.850000 365.000000 8.150000 ;
        RECT 360.000000 3.850000 365.000000 4.150000 ;
        RECT 410.000000 7.850000 415.000000 8.150000 ;
        RECT 410.000000 3.850000 415.000000 4.150000 ;
        RECT 460.000000 7.850000 465.000000 8.150000 ;
        RECT 460.000000 3.850000 465.000000 4.150000 ;
        RECT 510.000000 7.850000 515.000000 8.150000 ;
        RECT 510.000000 3.850000 515.000000 4.150000 ;
        RECT 560.000000 7.850000 565.000000 8.150000 ;
        RECT 560.000000 3.850000 565.000000 4.150000 ;
        RECT 18.000000 267.850000 28.000000 268.150000 ;
        RECT 18.000000 259.850000 28.000000 260.150000 ;
        RECT 18.000000 263.850000 28.000000 264.150000 ;
        RECT 60.000000 267.850000 65.000000 268.150000 ;
        RECT 60.000000 263.850000 65.000000 264.150000 ;
        RECT 60.000000 259.850000 65.000000 260.150000 ;
        RECT 110.000000 267.850000 115.000000 268.150000 ;
        RECT 110.000000 259.850000 115.000000 260.150000 ;
        RECT 110.000000 263.850000 115.000000 264.150000 ;
        RECT 18.000000 283.850000 28.000000 284.150000 ;
        RECT 18.000000 279.850000 28.000000 280.150000 ;
        RECT 18.000000 275.850000 28.000000 276.150000 ;
        RECT 18.000000 271.850000 28.000000 272.150000 ;
        RECT 18.000000 287.850000 28.000000 288.150000 ;
        RECT 18.000000 291.850000 28.000000 292.150000 ;
        RECT 18.000000 295.850000 28.000000 296.150000 ;
        RECT 18.000000 299.850000 28.000000 300.150000 ;
        RECT 18.000000 303.850000 28.000000 304.150000 ;
        RECT 60.000000 283.850000 65.000000 284.150000 ;
        RECT 60.000000 279.850000 65.000000 280.150000 ;
        RECT 60.000000 275.850000 65.000000 276.150000 ;
        RECT 60.000000 271.850000 65.000000 272.150000 ;
        RECT 60.000000 287.850000 65.000000 288.150000 ;
        RECT 60.000000 291.850000 65.000000 292.150000 ;
        RECT 60.000000 295.850000 65.000000 296.150000 ;
        RECT 60.000000 299.850000 65.000000 300.150000 ;
        RECT 60.000000 303.850000 65.000000 304.150000 ;
        RECT 18.000000 307.850000 28.000000 308.150000 ;
        RECT 18.000000 311.850000 28.000000 312.150000 ;
        RECT 18.000000 315.850000 28.000000 316.150000 ;
        RECT 18.000000 319.850000 28.000000 320.150000 ;
        RECT 18.000000 323.850000 28.000000 324.150000 ;
        RECT 18.000000 339.850000 28.000000 340.150000 ;
        RECT 18.000000 335.850000 28.000000 336.150000 ;
        RECT 18.000000 331.850000 28.000000 332.150000 ;
        RECT 18.000000 327.850000 28.000000 328.150000 ;
        RECT 60.000000 307.850000 65.000000 308.150000 ;
        RECT 60.000000 311.850000 65.000000 312.150000 ;
        RECT 60.000000 315.850000 65.000000 316.150000 ;
        RECT 60.000000 319.850000 65.000000 320.150000 ;
        RECT 60.000000 323.850000 65.000000 324.150000 ;
        RECT 60.000000 339.850000 65.000000 340.150000 ;
        RECT 60.000000 335.850000 65.000000 336.150000 ;
        RECT 60.000000 331.850000 65.000000 332.150000 ;
        RECT 60.000000 327.850000 65.000000 328.150000 ;
        RECT 110.000000 271.850000 115.000000 272.150000 ;
        RECT 110.000000 275.850000 115.000000 276.150000 ;
        RECT 110.000000 279.850000 115.000000 280.150000 ;
        RECT 110.000000 283.850000 115.000000 284.150000 ;
        RECT 110.000000 287.850000 115.000000 288.150000 ;
        RECT 110.000000 291.850000 115.000000 292.150000 ;
        RECT 110.000000 295.850000 115.000000 296.150000 ;
        RECT 110.000000 299.850000 115.000000 300.150000 ;
        RECT 110.000000 303.850000 115.000000 304.150000 ;
        RECT 110.000000 311.850000 115.000000 312.150000 ;
        RECT 110.000000 307.850000 115.000000 308.150000 ;
        RECT 110.000000 323.850000 115.000000 324.150000 ;
        RECT 110.000000 319.850000 115.000000 320.150000 ;
        RECT 110.000000 315.850000 115.000000 316.150000 ;
        RECT 110.000000 339.850000 115.000000 340.150000 ;
        RECT 110.000000 335.850000 115.000000 336.150000 ;
        RECT 110.000000 331.850000 115.000000 332.150000 ;
        RECT 110.000000 327.850000 115.000000 328.150000 ;
        RECT 160.000000 259.850000 165.000000 260.150000 ;
        RECT 160.000000 263.850000 165.000000 264.150000 ;
        RECT 160.000000 267.850000 165.000000 268.150000 ;
        RECT 210.000000 267.850000 215.000000 268.150000 ;
        RECT 210.000000 263.850000 215.000000 264.150000 ;
        RECT 210.000000 259.850000 215.000000 260.150000 ;
        RECT 260.000000 267.850000 265.000000 268.150000 ;
        RECT 260.000000 259.850000 265.000000 260.150000 ;
        RECT 260.000000 263.850000 265.000000 264.150000 ;
        RECT 160.000000 275.850000 165.000000 276.150000 ;
        RECT 160.000000 271.850000 165.000000 272.150000 ;
        RECT 160.000000 283.850000 165.000000 284.150000 ;
        RECT 160.000000 279.850000 165.000000 280.150000 ;
        RECT 160.000000 287.850000 165.000000 288.150000 ;
        RECT 160.000000 291.850000 165.000000 292.150000 ;
        RECT 160.000000 295.850000 165.000000 296.150000 ;
        RECT 160.000000 299.850000 165.000000 300.150000 ;
        RECT 160.000000 303.850000 165.000000 304.150000 ;
        RECT 210.000000 283.850000 215.000000 284.150000 ;
        RECT 210.000000 279.850000 215.000000 280.150000 ;
        RECT 210.000000 275.850000 215.000000 276.150000 ;
        RECT 210.000000 271.850000 215.000000 272.150000 ;
        RECT 210.000000 287.850000 215.000000 288.150000 ;
        RECT 210.000000 291.850000 215.000000 292.150000 ;
        RECT 210.000000 295.850000 215.000000 296.150000 ;
        RECT 210.000000 299.850000 215.000000 300.150000 ;
        RECT 210.000000 303.850000 215.000000 304.150000 ;
        RECT 160.000000 311.850000 165.000000 312.150000 ;
        RECT 160.000000 307.850000 165.000000 308.150000 ;
        RECT 160.000000 315.850000 165.000000 316.150000 ;
        RECT 160.000000 319.850000 165.000000 320.150000 ;
        RECT 160.000000 323.850000 165.000000 324.150000 ;
        RECT 160.000000 331.850000 165.000000 332.150000 ;
        RECT 160.000000 327.850000 165.000000 328.150000 ;
        RECT 160.000000 335.850000 165.000000 336.150000 ;
        RECT 160.000000 339.850000 165.000000 340.150000 ;
        RECT 210.000000 307.850000 215.000000 308.150000 ;
        RECT 210.000000 311.850000 215.000000 312.150000 ;
        RECT 210.000000 315.850000 215.000000 316.150000 ;
        RECT 210.000000 323.850000 215.000000 324.150000 ;
        RECT 210.000000 319.850000 215.000000 320.150000 ;
        RECT 210.000000 327.850000 215.000000 328.150000 ;
        RECT 210.000000 331.850000 215.000000 332.150000 ;
        RECT 210.000000 335.850000 215.000000 336.150000 ;
        RECT 210.000000 339.850000 215.000000 340.150000 ;
        RECT 260.000000 271.850000 265.000000 272.150000 ;
        RECT 260.000000 275.850000 265.000000 276.150000 ;
        RECT 260.000000 279.850000 265.000000 280.150000 ;
        RECT 260.000000 283.850000 265.000000 284.150000 ;
        RECT 260.000000 291.850000 265.000000 292.150000 ;
        RECT 260.000000 287.850000 265.000000 288.150000 ;
        RECT 260.000000 295.850000 265.000000 296.150000 ;
        RECT 260.000000 303.850000 265.000000 304.150000 ;
        RECT 260.000000 299.850000 265.000000 300.150000 ;
        RECT 260.000000 307.850000 265.000000 308.150000 ;
        RECT 260.000000 311.850000 265.000000 312.150000 ;
        RECT 260.000000 315.850000 265.000000 316.150000 ;
        RECT 260.000000 319.850000 265.000000 320.150000 ;
        RECT 260.000000 323.850000 265.000000 324.150000 ;
        RECT 260.000000 327.850000 265.000000 328.150000 ;
        RECT 260.000000 331.850000 265.000000 332.150000 ;
        RECT 260.000000 335.850000 265.000000 336.150000 ;
        RECT 260.000000 339.850000 265.000000 340.150000 ;
        RECT 310.000000 259.850000 315.000000 260.150000 ;
        RECT 310.000000 263.850000 315.000000 264.150000 ;
        RECT 310.000000 267.850000 315.000000 268.150000 ;
        RECT 360.000000 267.850000 365.000000 268.150000 ;
        RECT 360.000000 263.850000 365.000000 264.150000 ;
        RECT 360.000000 259.850000 365.000000 260.150000 ;
        RECT 410.000000 259.850000 415.000000 260.150000 ;
        RECT 410.000000 263.850000 415.000000 264.150000 ;
        RECT 410.000000 267.850000 415.000000 268.150000 ;
        RECT 310.000000 275.850000 315.000000 276.150000 ;
        RECT 310.000000 271.850000 315.000000 272.150000 ;
        RECT 310.000000 283.850000 315.000000 284.150000 ;
        RECT 310.000000 279.850000 315.000000 280.150000 ;
        RECT 310.000000 291.850000 315.000000 292.150000 ;
        RECT 310.000000 287.850000 315.000000 288.150000 ;
        RECT 310.000000 295.850000 315.000000 296.150000 ;
        RECT 310.000000 303.850000 315.000000 304.150000 ;
        RECT 310.000000 299.850000 315.000000 300.150000 ;
        RECT 360.000000 283.850000 365.000000 284.150000 ;
        RECT 360.000000 279.850000 365.000000 280.150000 ;
        RECT 360.000000 275.850000 365.000000 276.150000 ;
        RECT 360.000000 271.850000 365.000000 272.150000 ;
        RECT 360.000000 287.850000 365.000000 288.150000 ;
        RECT 360.000000 291.850000 365.000000 292.150000 ;
        RECT 360.000000 295.850000 365.000000 296.150000 ;
        RECT 360.000000 299.850000 365.000000 300.150000 ;
        RECT 360.000000 303.850000 365.000000 304.150000 ;
        RECT 310.000000 311.850000 315.000000 312.150000 ;
        RECT 310.000000 307.850000 315.000000 308.150000 ;
        RECT 310.000000 315.850000 315.000000 316.150000 ;
        RECT 310.000000 323.850000 315.000000 324.150000 ;
        RECT 310.000000 319.850000 315.000000 320.150000 ;
        RECT 310.000000 327.850000 315.000000 328.150000 ;
        RECT 310.000000 331.850000 315.000000 332.150000 ;
        RECT 310.000000 335.850000 315.000000 336.150000 ;
        RECT 310.000000 339.850000 315.000000 340.150000 ;
        RECT 360.000000 307.850000 365.000000 308.150000 ;
        RECT 360.000000 311.850000 365.000000 312.150000 ;
        RECT 360.000000 315.850000 365.000000 316.150000 ;
        RECT 360.000000 319.850000 365.000000 320.150000 ;
        RECT 360.000000 323.850000 365.000000 324.150000 ;
        RECT 360.000000 339.850000 365.000000 340.150000 ;
        RECT 360.000000 335.850000 365.000000 336.150000 ;
        RECT 360.000000 331.850000 365.000000 332.150000 ;
        RECT 360.000000 327.850000 365.000000 328.150000 ;
        RECT 410.000000 271.850000 415.000000 272.150000 ;
        RECT 410.000000 275.850000 415.000000 276.150000 ;
        RECT 410.000000 279.850000 415.000000 280.150000 ;
        RECT 410.000000 283.850000 415.000000 284.150000 ;
        RECT 410.000000 291.850000 415.000000 292.150000 ;
        RECT 410.000000 287.850000 415.000000 288.150000 ;
        RECT 410.000000 295.850000 415.000000 296.150000 ;
        RECT 410.000000 299.850000 415.000000 300.150000 ;
        RECT 410.000000 303.850000 415.000000 304.150000 ;
        RECT 410.000000 307.850000 415.000000 308.150000 ;
        RECT 410.000000 311.850000 415.000000 312.150000 ;
        RECT 410.000000 315.850000 415.000000 316.150000 ;
        RECT 410.000000 319.850000 415.000000 320.150000 ;
        RECT 410.000000 323.850000 415.000000 324.150000 ;
        RECT 410.000000 327.850000 415.000000 328.150000 ;
        RECT 410.000000 331.850000 415.000000 332.150000 ;
        RECT 410.000000 339.850000 415.000000 340.150000 ;
        RECT 410.000000 335.850000 415.000000 336.150000 ;
        RECT 460.000000 259.850000 465.000000 260.150000 ;
        RECT 460.000000 263.850000 465.000000 264.150000 ;
        RECT 460.000000 267.850000 465.000000 268.150000 ;
        RECT 510.000000 259.850000 515.000000 260.150000 ;
        RECT 510.000000 263.850000 515.000000 264.150000 ;
        RECT 510.000000 267.850000 515.000000 268.150000 ;
        RECT 560.000000 263.850000 565.000000 264.150000 ;
        RECT 560.000000 259.850000 565.000000 260.150000 ;
        RECT 560.000000 267.850000 565.000000 268.150000 ;
        RECT 460.000000 283.850000 465.000000 284.150000 ;
        RECT 460.000000 279.850000 465.000000 280.150000 ;
        RECT 460.000000 275.850000 465.000000 276.150000 ;
        RECT 460.000000 271.850000 465.000000 272.150000 ;
        RECT 460.000000 295.850000 465.000000 296.150000 ;
        RECT 460.000000 291.850000 465.000000 292.150000 ;
        RECT 460.000000 287.850000 465.000000 288.150000 ;
        RECT 510.000000 271.850000 515.000000 272.150000 ;
        RECT 510.000000 275.850000 515.000000 276.150000 ;
        RECT 510.000000 279.850000 515.000000 280.150000 ;
        RECT 510.000000 283.850000 515.000000 284.150000 ;
        RECT 510.000000 291.850000 515.000000 292.150000 ;
        RECT 510.000000 287.850000 515.000000 288.150000 ;
        RECT 510.000000 295.850000 515.000000 296.150000 ;
        RECT 510.000000 299.850000 515.000000 300.150000 ;
        RECT 510.000000 303.850000 515.000000 304.150000 ;
        RECT 460.000000 319.850000 465.000000 320.150000 ;
        RECT 460.000000 323.850000 465.000000 324.150000 ;
        RECT 460.000000 339.850000 465.000000 340.150000 ;
        RECT 460.000000 335.850000 465.000000 336.150000 ;
        RECT 460.000000 331.850000 465.000000 332.150000 ;
        RECT 460.000000 327.850000 465.000000 328.150000 ;
        RECT 510.000000 311.850000 515.000000 312.150000 ;
        RECT 510.000000 307.850000 515.000000 308.150000 ;
        RECT 510.000000 315.850000 515.000000 316.150000 ;
        RECT 510.000000 323.850000 515.000000 324.150000 ;
        RECT 510.000000 319.850000 515.000000 320.150000 ;
        RECT 510.000000 331.850000 515.000000 332.150000 ;
        RECT 510.000000 327.850000 515.000000 328.150000 ;
        RECT 510.000000 335.850000 515.000000 336.150000 ;
        RECT 510.000000 339.850000 515.000000 340.150000 ;
        RECT 560.000000 283.850000 565.000000 284.150000 ;
        RECT 560.000000 279.850000 565.000000 280.150000 ;
        RECT 560.000000 275.850000 565.000000 276.150000 ;
        RECT 560.000000 271.850000 565.000000 272.150000 ;
        RECT 560.000000 287.850000 565.000000 288.150000 ;
        RECT 560.000000 291.850000 565.000000 292.150000 ;
        RECT 560.000000 295.850000 565.000000 296.150000 ;
        RECT 560.000000 299.850000 565.000000 300.150000 ;
        RECT 560.000000 303.850000 565.000000 304.150000 ;
        RECT 560.000000 323.850000 565.000000 324.150000 ;
        RECT 560.000000 319.850000 565.000000 320.150000 ;
        RECT 560.000000 315.850000 565.000000 316.150000 ;
        RECT 560.000000 311.850000 565.000000 312.150000 ;
        RECT 560.000000 307.850000 565.000000 308.150000 ;
        RECT 560.000000 339.850000 565.000000 340.150000 ;
        RECT 560.000000 335.850000 565.000000 336.150000 ;
        RECT 560.000000 331.850000 565.000000 332.150000 ;
        RECT 560.000000 327.850000 565.000000 328.150000 ;
        RECT 610.000000 7.850000 615.000000 8.150000 ;
        RECT 610.000000 3.850000 615.000000 4.150000 ;
        RECT 660.000000 7.850000 665.000000 8.150000 ;
        RECT 660.000000 3.850000 665.000000 4.150000 ;
        RECT 710.000000 7.850000 715.000000 8.150000 ;
        RECT 710.000000 3.850000 715.000000 4.150000 ;
        RECT 760.000000 7.850000 765.000000 8.150000 ;
        RECT 760.000000 3.850000 765.000000 4.150000 ;
        RECT 810.000000 7.850000 815.000000 8.150000 ;
        RECT 810.000000 3.850000 815.000000 4.150000 ;
        RECT 860.000000 7.850000 865.000000 8.150000 ;
        RECT 860.000000 3.850000 865.000000 4.150000 ;
        RECT 960.000000 7.850000 965.000000 8.150000 ;
        RECT 960.000000 3.850000 965.000000 4.150000 ;
        RECT 910.000000 7.850000 915.000000 8.150000 ;
        RECT 910.000000 3.850000 915.000000 4.150000 ;
        RECT 1010.000000 7.850000 1015.000000 8.150000 ;
        RECT 1010.000000 3.850000 1015.000000 4.150000 ;
        RECT 1110.000000 7.850000 1115.000000 8.150000 ;
        RECT 1110.000000 3.850000 1115.000000 4.150000 ;
        RECT 1060.000000 7.850000 1065.000000 8.150000 ;
        RECT 1060.000000 3.850000 1065.000000 4.150000 ;
        RECT 1160.000000 3.850000 1165.000000 4.150000 ;
        RECT 1160.000000 7.850000 1165.000000 8.150000 ;
        RECT 1158.000000 27.850000 1168.000000 28.150000 ;
        RECT 1158.000000 23.850000 1168.000000 24.150000 ;
        RECT 1158.000000 19.850000 1168.000000 20.150000 ;
        RECT 1160.000000 15.850000 1165.000000 16.150000 ;
        RECT 1160.000000 11.850000 1165.000000 12.150000 ;
        RECT 1158.000000 31.850000 1168.000000 32.150000 ;
        RECT 1158.000000 35.850000 1168.000000 36.150000 ;
        RECT 1158.000000 43.850000 1168.000000 44.150000 ;
        RECT 1158.000000 39.850000 1168.000000 40.150000 ;
        RECT 610.000000 267.850000 615.000000 268.150000 ;
        RECT 610.000000 263.850000 615.000000 264.150000 ;
        RECT 610.000000 259.850000 615.000000 260.150000 ;
        RECT 660.000000 259.850000 665.000000 260.150000 ;
        RECT 660.000000 263.850000 665.000000 264.150000 ;
        RECT 660.000000 267.850000 665.000000 268.150000 ;
        RECT 710.000000 267.850000 715.000000 268.150000 ;
        RECT 710.000000 259.850000 715.000000 260.150000 ;
        RECT 710.000000 263.850000 715.000000 264.150000 ;
        RECT 610.000000 283.850000 615.000000 284.150000 ;
        RECT 610.000000 279.850000 615.000000 280.150000 ;
        RECT 610.000000 275.850000 615.000000 276.150000 ;
        RECT 610.000000 271.850000 615.000000 272.150000 ;
        RECT 610.000000 287.850000 615.000000 288.150000 ;
        RECT 610.000000 291.850000 615.000000 292.150000 ;
        RECT 610.000000 295.850000 615.000000 296.150000 ;
        RECT 610.000000 299.850000 615.000000 300.150000 ;
        RECT 610.000000 303.850000 615.000000 304.150000 ;
        RECT 660.000000 275.850000 665.000000 276.150000 ;
        RECT 660.000000 271.850000 665.000000 272.150000 ;
        RECT 660.000000 283.850000 665.000000 284.150000 ;
        RECT 660.000000 279.850000 665.000000 280.150000 ;
        RECT 660.000000 287.850000 665.000000 288.150000 ;
        RECT 660.000000 291.850000 665.000000 292.150000 ;
        RECT 660.000000 295.850000 665.000000 296.150000 ;
        RECT 660.000000 303.850000 665.000000 304.150000 ;
        RECT 660.000000 299.850000 665.000000 300.150000 ;
        RECT 610.000000 307.850000 615.000000 308.150000 ;
        RECT 610.000000 311.850000 615.000000 312.150000 ;
        RECT 610.000000 315.850000 615.000000 316.150000 ;
        RECT 610.000000 319.850000 615.000000 320.150000 ;
        RECT 610.000000 323.850000 615.000000 324.150000 ;
        RECT 610.000000 339.850000 615.000000 340.150000 ;
        RECT 610.000000 335.850000 615.000000 336.150000 ;
        RECT 610.000000 331.850000 615.000000 332.150000 ;
        RECT 610.000000 327.850000 615.000000 328.150000 ;
        RECT 660.000000 311.850000 665.000000 312.150000 ;
        RECT 660.000000 307.850000 665.000000 308.150000 ;
        RECT 660.000000 315.850000 665.000000 316.150000 ;
        RECT 660.000000 319.850000 665.000000 320.150000 ;
        RECT 660.000000 323.850000 665.000000 324.150000 ;
        RECT 660.000000 331.850000 665.000000 332.150000 ;
        RECT 660.000000 327.850000 665.000000 328.150000 ;
        RECT 660.000000 335.850000 665.000000 336.150000 ;
        RECT 660.000000 339.850000 665.000000 340.150000 ;
        RECT 710.000000 271.850000 715.000000 272.150000 ;
        RECT 710.000000 275.850000 715.000000 276.150000 ;
        RECT 710.000000 279.850000 715.000000 280.150000 ;
        RECT 710.000000 283.850000 715.000000 284.150000 ;
        RECT 710.000000 287.850000 715.000000 288.150000 ;
        RECT 710.000000 291.850000 715.000000 292.150000 ;
        RECT 710.000000 295.850000 715.000000 296.150000 ;
        RECT 710.000000 299.850000 715.000000 300.150000 ;
        RECT 710.000000 303.850000 715.000000 304.150000 ;
        RECT 710.000000 323.850000 715.000000 324.150000 ;
        RECT 710.000000 319.850000 715.000000 320.150000 ;
        RECT 710.000000 315.850000 715.000000 316.150000 ;
        RECT 710.000000 311.850000 715.000000 312.150000 ;
        RECT 710.000000 307.850000 715.000000 308.150000 ;
        RECT 710.000000 339.850000 715.000000 340.150000 ;
        RECT 710.000000 335.850000 715.000000 336.150000 ;
        RECT 710.000000 331.850000 715.000000 332.150000 ;
        RECT 710.000000 327.850000 715.000000 328.150000 ;
        RECT 760.000000 267.850000 765.000000 268.150000 ;
        RECT 760.000000 263.850000 765.000000 264.150000 ;
        RECT 760.000000 259.850000 765.000000 260.150000 ;
        RECT 810.000000 259.850000 815.000000 260.150000 ;
        RECT 810.000000 263.850000 815.000000 264.150000 ;
        RECT 810.000000 267.850000 815.000000 268.150000 ;
        RECT 860.000000 267.850000 865.000000 268.150000 ;
        RECT 860.000000 259.850000 865.000000 260.150000 ;
        RECT 860.000000 263.850000 865.000000 264.150000 ;
        RECT 760.000000 283.850000 765.000000 284.150000 ;
        RECT 760.000000 279.850000 765.000000 280.150000 ;
        RECT 760.000000 275.850000 765.000000 276.150000 ;
        RECT 760.000000 271.850000 765.000000 272.150000 ;
        RECT 760.000000 287.850000 765.000000 288.150000 ;
        RECT 760.000000 291.850000 765.000000 292.150000 ;
        RECT 760.000000 295.850000 765.000000 296.150000 ;
        RECT 760.000000 299.850000 765.000000 300.150000 ;
        RECT 760.000000 303.850000 765.000000 304.150000 ;
        RECT 810.000000 275.850000 815.000000 276.150000 ;
        RECT 810.000000 271.850000 815.000000 272.150000 ;
        RECT 810.000000 283.850000 815.000000 284.150000 ;
        RECT 810.000000 279.850000 815.000000 280.150000 ;
        RECT 810.000000 287.850000 815.000000 288.150000 ;
        RECT 810.000000 291.850000 815.000000 292.150000 ;
        RECT 810.000000 295.850000 815.000000 296.150000 ;
        RECT 810.000000 303.850000 815.000000 304.150000 ;
        RECT 810.000000 299.850000 815.000000 300.150000 ;
        RECT 760.000000 307.850000 765.000000 308.150000 ;
        RECT 760.000000 311.850000 765.000000 312.150000 ;
        RECT 760.000000 315.850000 765.000000 316.150000 ;
        RECT 760.000000 319.850000 765.000000 320.150000 ;
        RECT 760.000000 323.850000 765.000000 324.150000 ;
        RECT 760.000000 339.850000 765.000000 340.150000 ;
        RECT 760.000000 335.850000 765.000000 336.150000 ;
        RECT 760.000000 331.850000 765.000000 332.150000 ;
        RECT 760.000000 327.850000 765.000000 328.150000 ;
        RECT 810.000000 311.850000 815.000000 312.150000 ;
        RECT 810.000000 307.850000 815.000000 308.150000 ;
        RECT 810.000000 315.850000 815.000000 316.150000 ;
        RECT 810.000000 319.850000 815.000000 320.150000 ;
        RECT 810.000000 323.850000 815.000000 324.150000 ;
        RECT 810.000000 331.850000 815.000000 332.150000 ;
        RECT 810.000000 327.850000 815.000000 328.150000 ;
        RECT 810.000000 335.850000 815.000000 336.150000 ;
        RECT 810.000000 339.850000 815.000000 340.150000 ;
        RECT 860.000000 271.850000 865.000000 272.150000 ;
        RECT 860.000000 275.850000 865.000000 276.150000 ;
        RECT 860.000000 279.850000 865.000000 280.150000 ;
        RECT 860.000000 283.850000 865.000000 284.150000 ;
        RECT 860.000000 287.850000 865.000000 288.150000 ;
        RECT 860.000000 291.850000 865.000000 292.150000 ;
        RECT 860.000000 295.850000 865.000000 296.150000 ;
        RECT 860.000000 299.850000 865.000000 300.150000 ;
        RECT 860.000000 303.850000 865.000000 304.150000 ;
        RECT 860.000000 323.850000 865.000000 324.150000 ;
        RECT 860.000000 319.850000 865.000000 320.150000 ;
        RECT 860.000000 315.850000 865.000000 316.150000 ;
        RECT 860.000000 311.850000 865.000000 312.150000 ;
        RECT 860.000000 307.850000 865.000000 308.150000 ;
        RECT 860.000000 339.850000 865.000000 340.150000 ;
        RECT 860.000000 335.850000 865.000000 336.150000 ;
        RECT 860.000000 331.850000 865.000000 332.150000 ;
        RECT 860.000000 327.850000 865.000000 328.150000 ;
        RECT 1158.000000 47.850000 1168.000000 48.150000 ;
        RECT 1158.000000 51.850000 1168.000000 52.150000 ;
        RECT 1158.000000 63.850000 1168.000000 64.150000 ;
        RECT 1158.000000 59.850000 1168.000000 60.150000 ;
        RECT 1158.000000 55.850000 1168.000000 56.150000 ;
        RECT 1158.000000 67.850000 1168.000000 68.150000 ;
        RECT 1158.000000 71.850000 1168.000000 72.150000 ;
        RECT 1158.000000 79.850000 1168.000000 80.150000 ;
        RECT 1158.000000 75.850000 1168.000000 76.150000 ;
        RECT 1158.000000 83.850000 1168.000000 84.150000 ;
        RECT 1158.000000 87.850000 1168.000000 88.150000 ;
        RECT 1158.000000 91.850000 1168.000000 92.150000 ;
        RECT 1158.000000 99.850000 1168.000000 100.150000 ;
        RECT 1158.000000 95.850000 1168.000000 96.150000 ;
        RECT 1158.000000 103.850000 1168.000000 104.150000 ;
        RECT 1158.000000 107.850000 1168.000000 108.150000 ;
        RECT 1158.000000 119.850000 1168.000000 120.150000 ;
        RECT 1158.000000 115.850000 1168.000000 116.150000 ;
        RECT 1158.000000 111.850000 1168.000000 112.150000 ;
        RECT 1158.000000 123.850000 1168.000000 124.150000 ;
        RECT 1158.000000 127.850000 1168.000000 128.150000 ;
        RECT 1158.000000 135.850000 1168.000000 136.150000 ;
        RECT 1158.000000 131.850000 1168.000000 132.150000 ;
        RECT 1158.000000 139.850000 1168.000000 140.150000 ;
        RECT 1158.000000 143.850000 1168.000000 144.150000 ;
        RECT 1158.000000 147.850000 1168.000000 148.150000 ;
        RECT 1158.000000 155.850000 1168.000000 156.150000 ;
        RECT 1158.000000 151.850000 1168.000000 152.150000 ;
        RECT 1158.000000 159.850000 1168.000000 160.150000 ;
        RECT 1158.000000 163.850000 1168.000000 164.150000 ;
        RECT 1158.000000 175.850000 1168.000000 176.150000 ;
        RECT 1158.000000 171.850000 1168.000000 172.150000 ;
        RECT 1158.000000 167.850000 1168.000000 168.150000 ;
        RECT 1158.000000 179.850000 1168.000000 180.150000 ;
        RECT 1158.000000 183.850000 1168.000000 184.150000 ;
        RECT 1158.000000 191.850000 1168.000000 192.150000 ;
        RECT 1158.000000 187.850000 1168.000000 188.150000 ;
        RECT 960.000000 267.850000 965.000000 268.150000 ;
        RECT 960.000000 263.850000 965.000000 264.150000 ;
        RECT 960.000000 259.850000 965.000000 260.150000 ;
        RECT 910.000000 267.850000 915.000000 268.150000 ;
        RECT 910.000000 263.850000 915.000000 264.150000 ;
        RECT 910.000000 259.850000 915.000000 260.150000 ;
        RECT 1010.000000 259.850000 1015.000000 260.150000 ;
        RECT 1010.000000 263.850000 1015.000000 264.150000 ;
        RECT 1010.000000 267.850000 1015.000000 268.150000 ;
        RECT 960.000000 283.850000 965.000000 284.150000 ;
        RECT 960.000000 279.850000 965.000000 280.150000 ;
        RECT 960.000000 275.850000 965.000000 276.150000 ;
        RECT 960.000000 271.850000 965.000000 272.150000 ;
        RECT 960.000000 287.850000 965.000000 288.150000 ;
        RECT 960.000000 291.850000 965.000000 292.150000 ;
        RECT 960.000000 295.850000 965.000000 296.150000 ;
        RECT 960.000000 299.850000 965.000000 300.150000 ;
        RECT 960.000000 303.850000 965.000000 304.150000 ;
        RECT 960.000000 311.850000 965.000000 312.150000 ;
        RECT 960.000000 307.850000 965.000000 308.150000 ;
        RECT 960.000000 323.850000 965.000000 324.150000 ;
        RECT 960.000000 319.850000 965.000000 320.150000 ;
        RECT 960.000000 315.850000 965.000000 316.150000 ;
        RECT 960.000000 339.850000 965.000000 340.150000 ;
        RECT 960.000000 335.850000 965.000000 336.150000 ;
        RECT 960.000000 331.850000 965.000000 332.150000 ;
        RECT 960.000000 327.850000 965.000000 328.150000 ;
        RECT 910.000000 283.850000 915.000000 284.150000 ;
        RECT 910.000000 279.850000 915.000000 280.150000 ;
        RECT 910.000000 275.850000 915.000000 276.150000 ;
        RECT 910.000000 271.850000 915.000000 272.150000 ;
        RECT 910.000000 287.850000 915.000000 288.150000 ;
        RECT 910.000000 291.850000 915.000000 292.150000 ;
        RECT 910.000000 295.850000 915.000000 296.150000 ;
        RECT 910.000000 299.850000 915.000000 300.150000 ;
        RECT 910.000000 303.850000 915.000000 304.150000 ;
        RECT 910.000000 307.850000 915.000000 308.150000 ;
        RECT 910.000000 311.850000 915.000000 312.150000 ;
        RECT 910.000000 315.850000 915.000000 316.150000 ;
        RECT 910.000000 319.850000 915.000000 320.150000 ;
        RECT 910.000000 323.850000 915.000000 324.150000 ;
        RECT 910.000000 339.850000 915.000000 340.150000 ;
        RECT 910.000000 335.850000 915.000000 336.150000 ;
        RECT 910.000000 331.850000 915.000000 332.150000 ;
        RECT 910.000000 327.850000 915.000000 328.150000 ;
        RECT 1010.000000 275.850000 1015.000000 276.150000 ;
        RECT 1010.000000 271.850000 1015.000000 272.150000 ;
        RECT 1010.000000 283.850000 1015.000000 284.150000 ;
        RECT 1010.000000 279.850000 1015.000000 280.150000 ;
        RECT 1010.000000 287.850000 1015.000000 288.150000 ;
        RECT 1010.000000 291.850000 1015.000000 292.150000 ;
        RECT 1010.000000 295.850000 1015.000000 296.150000 ;
        RECT 1010.000000 303.850000 1015.000000 304.150000 ;
        RECT 1010.000000 299.850000 1015.000000 300.150000 ;
        RECT 1010.000000 311.850000 1015.000000 312.150000 ;
        RECT 1010.000000 307.850000 1015.000000 308.150000 ;
        RECT 1010.000000 315.850000 1015.000000 316.150000 ;
        RECT 1010.000000 319.850000 1015.000000 320.150000 ;
        RECT 1010.000000 323.850000 1015.000000 324.150000 ;
        RECT 1010.000000 331.850000 1015.000000 332.150000 ;
        RECT 1010.000000 327.850000 1015.000000 328.150000 ;
        RECT 1010.000000 335.850000 1015.000000 336.150000 ;
        RECT 1010.000000 339.850000 1015.000000 340.150000 ;
        RECT 1110.000000 267.850000 1115.000000 268.150000 ;
        RECT 1110.000000 263.850000 1115.000000 264.150000 ;
        RECT 1110.000000 259.850000 1115.000000 260.150000 ;
        RECT 1060.000000 267.850000 1065.000000 268.150000 ;
        RECT 1060.000000 263.850000 1065.000000 264.150000 ;
        RECT 1060.000000 259.850000 1065.000000 260.150000 ;
        RECT 1158.000000 203.850000 1168.000000 204.150000 ;
        RECT 1158.000000 195.850000 1168.000000 196.150000 ;
        RECT 1158.000000 199.850000 1168.000000 200.150000 ;
        RECT 1158.000000 211.850000 1168.000000 212.150000 ;
        RECT 1158.000000 207.850000 1168.000000 208.150000 ;
        RECT 1158.000000 215.850000 1168.000000 216.150000 ;
        RECT 1158.000000 219.850000 1168.000000 220.150000 ;
        RECT 1158.000000 227.850000 1168.000000 228.150000 ;
        RECT 1158.000000 223.850000 1168.000000 224.150000 ;
        RECT 1158.000000 231.850000 1168.000000 232.150000 ;
        RECT 1158.000000 235.850000 1168.000000 236.150000 ;
        RECT 1158.000000 239.850000 1168.000000 240.150000 ;
        RECT 1158.000000 247.850000 1168.000000 248.150000 ;
        RECT 1158.000000 243.850000 1168.000000 244.150000 ;
        RECT 1158.000000 251.850000 1168.000000 252.150000 ;
        RECT 1158.000000 255.850000 1168.000000 256.150000 ;
        RECT 1158.000000 267.850000 1168.000000 268.150000 ;
        RECT 1158.000000 259.850000 1168.000000 260.150000 ;
        RECT 1158.000000 263.850000 1168.000000 264.150000 ;
        RECT 1110.000000 283.850000 1115.000000 284.150000 ;
        RECT 1110.000000 279.850000 1115.000000 280.150000 ;
        RECT 1110.000000 275.850000 1115.000000 276.150000 ;
        RECT 1110.000000 271.850000 1115.000000 272.150000 ;
        RECT 1110.000000 287.850000 1115.000000 288.150000 ;
        RECT 1110.000000 291.850000 1115.000000 292.150000 ;
        RECT 1110.000000 295.850000 1115.000000 296.150000 ;
        RECT 1110.000000 299.850000 1115.000000 300.150000 ;
        RECT 1110.000000 303.850000 1115.000000 304.150000 ;
        RECT 1110.000000 311.850000 1115.000000 312.150000 ;
        RECT 1110.000000 307.850000 1115.000000 308.150000 ;
        RECT 1110.000000 323.850000 1115.000000 324.150000 ;
        RECT 1110.000000 319.850000 1115.000000 320.150000 ;
        RECT 1110.000000 315.850000 1115.000000 316.150000 ;
        RECT 1110.000000 339.850000 1115.000000 340.150000 ;
        RECT 1110.000000 335.850000 1115.000000 336.150000 ;
        RECT 1110.000000 331.850000 1115.000000 332.150000 ;
        RECT 1110.000000 327.850000 1115.000000 328.150000 ;
        RECT 1060.000000 283.850000 1065.000000 284.150000 ;
        RECT 1060.000000 279.850000 1065.000000 280.150000 ;
        RECT 1060.000000 275.850000 1065.000000 276.150000 ;
        RECT 1060.000000 271.850000 1065.000000 272.150000 ;
        RECT 1060.000000 287.850000 1065.000000 288.150000 ;
        RECT 1060.000000 291.850000 1065.000000 292.150000 ;
        RECT 1060.000000 295.850000 1065.000000 296.150000 ;
        RECT 1060.000000 299.850000 1065.000000 300.150000 ;
        RECT 1060.000000 303.850000 1065.000000 304.150000 ;
        RECT 1060.000000 307.850000 1065.000000 308.150000 ;
        RECT 1060.000000 311.850000 1065.000000 312.150000 ;
        RECT 1060.000000 315.850000 1065.000000 316.150000 ;
        RECT 1060.000000 319.850000 1065.000000 320.150000 ;
        RECT 1060.000000 323.850000 1065.000000 324.150000 ;
        RECT 1060.000000 339.850000 1065.000000 340.150000 ;
        RECT 1060.000000 335.850000 1065.000000 336.150000 ;
        RECT 1060.000000 331.850000 1065.000000 332.150000 ;
        RECT 1060.000000 327.850000 1065.000000 328.150000 ;
        RECT 1158.000000 283.850000 1168.000000 284.150000 ;
        RECT 1158.000000 279.850000 1168.000000 280.150000 ;
        RECT 1158.000000 275.850000 1168.000000 276.150000 ;
        RECT 1158.000000 271.850000 1168.000000 272.150000 ;
        RECT 1158.000000 287.850000 1168.000000 288.150000 ;
        RECT 1158.000000 291.850000 1168.000000 292.150000 ;
        RECT 1158.000000 295.850000 1168.000000 296.150000 ;
        RECT 1158.000000 299.850000 1168.000000 300.150000 ;
        RECT 1158.000000 303.850000 1168.000000 304.150000 ;
        RECT 1158.000000 307.850000 1168.000000 308.150000 ;
        RECT 1158.000000 311.850000 1168.000000 312.150000 ;
        RECT 1158.000000 315.850000 1168.000000 316.150000 ;
        RECT 1158.000000 319.850000 1168.000000 320.150000 ;
        RECT 1158.000000 323.850000 1168.000000 324.150000 ;
        RECT 1158.000000 339.850000 1168.000000 340.150000 ;
        RECT 1158.000000 335.850000 1168.000000 336.150000 ;
        RECT 1158.000000 331.850000 1168.000000 332.150000 ;
        RECT 1158.000000 327.850000 1168.000000 328.150000 ;
        RECT 60.000000 379.850000 65.000000 380.150000 ;
        RECT 18.000000 379.850000 28.000000 380.150000 ;
        RECT 18.000000 343.850000 28.000000 344.150000 ;
        RECT 18.000000 347.850000 28.000000 348.150000 ;
        RECT 18.000000 351.850000 28.000000 352.150000 ;
        RECT 18.000000 359.850000 28.000000 360.150000 ;
        RECT 18.000000 355.850000 28.000000 356.150000 ;
        RECT 18.000000 375.850000 28.000000 376.150000 ;
        RECT 18.000000 371.850000 28.000000 372.150000 ;
        RECT 18.000000 367.850000 28.000000 368.150000 ;
        RECT 18.000000 363.850000 28.000000 364.150000 ;
        RECT 60.000000 347.850000 65.000000 348.150000 ;
        RECT 60.000000 343.850000 65.000000 344.150000 ;
        RECT 60.000000 375.850000 65.000000 376.150000 ;
        RECT 60.000000 371.850000 65.000000 372.150000 ;
        RECT 60.000000 367.850000 65.000000 368.150000 ;
        RECT 60.000000 363.850000 65.000000 364.150000 ;
        RECT 18.000000 395.850000 28.000000 396.150000 ;
        RECT 18.000000 391.850000 28.000000 392.150000 ;
        RECT 18.000000 387.850000 28.000000 388.150000 ;
        RECT 18.000000 383.850000 28.000000 384.150000 ;
        RECT 18.000000 407.850000 28.000000 408.150000 ;
        RECT 18.000000 399.850000 28.000000 400.150000 ;
        RECT 18.000000 403.850000 28.000000 404.150000 ;
        RECT 18.000000 411.850000 28.000000 412.150000 ;
        RECT 18.000000 415.850000 28.000000 416.150000 ;
        RECT 60.000000 395.850000 65.000000 396.150000 ;
        RECT 60.000000 391.850000 65.000000 392.150000 ;
        RECT 60.000000 387.850000 65.000000 388.150000 ;
        RECT 60.000000 383.850000 65.000000 384.150000 ;
        RECT 60.000000 407.850000 65.000000 408.150000 ;
        RECT 60.000000 399.850000 65.000000 400.150000 ;
        RECT 60.000000 403.850000 65.000000 404.150000 ;
        RECT 60.000000 411.850000 65.000000 412.150000 ;
        RECT 60.000000 415.850000 65.000000 416.150000 ;
        RECT 110.000000 379.850000 115.000000 380.150000 ;
        RECT 110.000000 351.850000 115.000000 352.150000 ;
        RECT 110.000000 347.850000 115.000000 348.150000 ;
        RECT 110.000000 343.850000 115.000000 344.150000 ;
        RECT 110.000000 359.850000 115.000000 360.150000 ;
        RECT 110.000000 355.850000 115.000000 356.150000 ;
        RECT 110.000000 375.850000 115.000000 376.150000 ;
        RECT 110.000000 371.850000 115.000000 372.150000 ;
        RECT 110.000000 367.850000 115.000000 368.150000 ;
        RECT 110.000000 363.850000 115.000000 364.150000 ;
        RECT 110.000000 383.850000 115.000000 384.150000 ;
        RECT 110.000000 387.850000 115.000000 388.150000 ;
        RECT 110.000000 391.850000 115.000000 392.150000 ;
        RECT 110.000000 395.850000 115.000000 396.150000 ;
        RECT 110.000000 407.850000 115.000000 408.150000 ;
        RECT 110.000000 399.850000 115.000000 400.150000 ;
        RECT 110.000000 403.850000 115.000000 404.150000 ;
        RECT 110.000000 411.850000 115.000000 412.150000 ;
        RECT 110.000000 415.850000 115.000000 416.150000 ;
        RECT 18.000000 431.850000 28.000000 432.150000 ;
        RECT 18.000000 427.850000 28.000000 428.150000 ;
        RECT 18.000000 423.850000 28.000000 424.150000 ;
        RECT 18.000000 419.850000 28.000000 420.150000 ;
        RECT 18.000000 435.850000 28.000000 436.150000 ;
        RECT 18.000000 439.850000 28.000000 440.150000 ;
        RECT 18.000000 443.850000 28.000000 444.150000 ;
        RECT 18.000000 447.850000 28.000000 448.150000 ;
        RECT 18.000000 451.850000 28.000000 452.150000 ;
        RECT 60.000000 431.850000 65.000000 432.150000 ;
        RECT 60.000000 427.850000 65.000000 428.150000 ;
        RECT 60.000000 423.850000 65.000000 424.150000 ;
        RECT 60.000000 419.850000 65.000000 420.150000 ;
        RECT 60.000000 435.850000 65.000000 436.150000 ;
        RECT 60.000000 439.850000 65.000000 440.150000 ;
        RECT 60.000000 443.850000 65.000000 444.150000 ;
        RECT 60.000000 447.850000 65.000000 448.150000 ;
        RECT 60.000000 451.850000 65.000000 452.150000 ;
        RECT 18.000000 455.850000 28.000000 456.150000 ;
        RECT 18.000000 459.850000 28.000000 460.150000 ;
        RECT 18.000000 463.850000 28.000000 464.150000 ;
        RECT 18.000000 467.850000 28.000000 468.150000 ;
        RECT 18.000000 471.850000 28.000000 472.150000 ;
        RECT 18.000000 487.850000 28.000000 488.150000 ;
        RECT 18.000000 483.850000 28.000000 484.150000 ;
        RECT 18.000000 479.850000 28.000000 480.150000 ;
        RECT 18.000000 475.850000 28.000000 476.150000 ;
        RECT 60.000000 455.850000 65.000000 456.150000 ;
        RECT 60.000000 459.850000 65.000000 460.150000 ;
        RECT 60.000000 463.850000 65.000000 464.150000 ;
        RECT 60.000000 467.850000 65.000000 468.150000 ;
        RECT 60.000000 471.850000 65.000000 472.150000 ;
        RECT 60.000000 487.850000 65.000000 488.150000 ;
        RECT 60.000000 483.850000 65.000000 484.150000 ;
        RECT 60.000000 479.850000 65.000000 480.150000 ;
        RECT 60.000000 475.850000 65.000000 476.150000 ;
        RECT 110.000000 419.850000 115.000000 420.150000 ;
        RECT 110.000000 423.850000 115.000000 424.150000 ;
        RECT 110.000000 427.850000 115.000000 428.150000 ;
        RECT 110.000000 431.850000 115.000000 432.150000 ;
        RECT 110.000000 435.850000 115.000000 436.150000 ;
        RECT 110.000000 439.850000 115.000000 440.150000 ;
        RECT 110.000000 443.850000 115.000000 444.150000 ;
        RECT 110.000000 447.850000 115.000000 448.150000 ;
        RECT 110.000000 451.850000 115.000000 452.150000 ;
        RECT 110.000000 459.850000 115.000000 460.150000 ;
        RECT 110.000000 455.850000 115.000000 456.150000 ;
        RECT 110.000000 471.850000 115.000000 472.150000 ;
        RECT 110.000000 467.850000 115.000000 468.150000 ;
        RECT 110.000000 463.850000 115.000000 464.150000 ;
        RECT 110.000000 487.850000 115.000000 488.150000 ;
        RECT 110.000000 483.850000 115.000000 484.150000 ;
        RECT 110.000000 479.850000 115.000000 480.150000 ;
        RECT 110.000000 475.850000 115.000000 476.150000 ;
        RECT 210.000000 379.850000 215.000000 380.150000 ;
        RECT 160.000000 379.850000 165.000000 380.150000 ;
        RECT 160.000000 343.850000 165.000000 344.150000 ;
        RECT 160.000000 347.850000 165.000000 348.150000 ;
        RECT 160.000000 351.850000 165.000000 352.150000 ;
        RECT 160.000000 359.850000 165.000000 360.150000 ;
        RECT 160.000000 355.850000 165.000000 356.150000 ;
        RECT 160.000000 363.850000 165.000000 364.150000 ;
        RECT 160.000000 367.850000 165.000000 368.150000 ;
        RECT 160.000000 371.850000 165.000000 372.150000 ;
        RECT 160.000000 375.850000 165.000000 376.150000 ;
        RECT 210.000000 343.850000 215.000000 344.150000 ;
        RECT 210.000000 347.850000 215.000000 348.150000 ;
        RECT 210.000000 351.850000 215.000000 352.150000 ;
        RECT 210.000000 355.850000 215.000000 356.150000 ;
        RECT 210.000000 359.850000 215.000000 360.150000 ;
        RECT 210.000000 375.850000 215.000000 376.150000 ;
        RECT 210.000000 371.850000 215.000000 372.150000 ;
        RECT 210.000000 367.850000 215.000000 368.150000 ;
        RECT 210.000000 363.850000 215.000000 364.150000 ;
        RECT 160.000000 387.850000 165.000000 388.150000 ;
        RECT 160.000000 383.850000 165.000000 384.150000 ;
        RECT 160.000000 391.850000 165.000000 392.150000 ;
        RECT 160.000000 395.850000 165.000000 396.150000 ;
        RECT 160.000000 399.850000 165.000000 400.150000 ;
        RECT 210.000000 383.850000 215.000000 384.150000 ;
        RECT 210.000000 387.850000 215.000000 388.150000 ;
        RECT 210.000000 391.850000 215.000000 392.150000 ;
        RECT 210.000000 395.850000 215.000000 396.150000 ;
        RECT 210.000000 407.850000 215.000000 408.150000 ;
        RECT 210.000000 399.850000 215.000000 400.150000 ;
        RECT 210.000000 403.850000 215.000000 404.150000 ;
        RECT 210.000000 411.850000 215.000000 412.150000 ;
        RECT 210.000000 415.850000 215.000000 416.150000 ;
        RECT 260.000000 379.850000 265.000000 380.150000 ;
        RECT 260.000000 343.850000 265.000000 344.150000 ;
        RECT 260.000000 347.850000 265.000000 348.150000 ;
        RECT 260.000000 351.850000 265.000000 352.150000 ;
        RECT 260.000000 355.850000 265.000000 356.150000 ;
        RECT 260.000000 359.850000 265.000000 360.150000 ;
        RECT 260.000000 363.850000 265.000000 364.150000 ;
        RECT 260.000000 367.850000 265.000000 368.150000 ;
        RECT 260.000000 371.850000 265.000000 372.150000 ;
        RECT 260.000000 375.850000 265.000000 376.150000 ;
        RECT 260.000000 383.850000 265.000000 384.150000 ;
        RECT 260.000000 387.850000 265.000000 388.150000 ;
        RECT 260.000000 391.850000 265.000000 392.150000 ;
        RECT 260.000000 395.850000 265.000000 396.150000 ;
        RECT 260.000000 399.850000 265.000000 400.150000 ;
        RECT 210.000000 431.850000 215.000000 432.150000 ;
        RECT 210.000000 427.850000 215.000000 428.150000 ;
        RECT 210.000000 423.850000 215.000000 424.150000 ;
        RECT 210.000000 419.850000 215.000000 420.150000 ;
        RECT 210.000000 435.850000 215.000000 436.150000 ;
        RECT 210.000000 439.850000 215.000000 440.150000 ;
        RECT 210.000000 443.850000 215.000000 444.150000 ;
        RECT 210.000000 447.850000 215.000000 448.150000 ;
        RECT 210.000000 451.850000 215.000000 452.150000 ;
        RECT 160.000000 463.850000 165.000000 464.150000 ;
        RECT 160.000000 467.850000 165.000000 468.150000 ;
        RECT 160.000000 471.850000 165.000000 472.150000 ;
        RECT 160.000000 479.850000 165.000000 480.150000 ;
        RECT 160.000000 475.850000 165.000000 476.150000 ;
        RECT 160.000000 487.850000 165.000000 488.150000 ;
        RECT 160.000000 483.850000 165.000000 484.150000 ;
        RECT 210.000000 455.850000 215.000000 456.150000 ;
        RECT 210.000000 459.850000 215.000000 460.150000 ;
        RECT 210.000000 463.850000 215.000000 464.150000 ;
        RECT 210.000000 467.850000 215.000000 468.150000 ;
        RECT 210.000000 471.850000 215.000000 472.150000 ;
        RECT 210.000000 475.850000 215.000000 476.150000 ;
        RECT 210.000000 479.850000 215.000000 480.150000 ;
        RECT 210.000000 483.850000 215.000000 484.150000 ;
        RECT 210.000000 487.850000 215.000000 488.150000 ;
        RECT 260.000000 467.850000 265.000000 468.150000 ;
        RECT 260.000000 463.850000 265.000000 464.150000 ;
        RECT 260.000000 471.850000 265.000000 472.150000 ;
        RECT 260.000000 475.850000 265.000000 476.150000 ;
        RECT 260.000000 479.850000 265.000000 480.150000 ;
        RECT 260.000000 487.850000 265.000000 488.150000 ;
        RECT 260.000000 483.850000 265.000000 484.150000 ;
        RECT 18.000000 491.850000 28.000000 492.150000 ;
        RECT 18.000000 495.850000 28.000000 496.150000 ;
        RECT 18.000000 499.850000 28.000000 500.150000 ;
        RECT 18.000000 503.850000 28.000000 504.150000 ;
        RECT 18.000000 507.850000 28.000000 508.150000 ;
        RECT 18.000000 515.850000 28.000000 516.150000 ;
        RECT 18.000000 511.850000 28.000000 512.150000 ;
        RECT 60.000000 491.850000 65.000000 492.150000 ;
        RECT 60.000000 495.850000 65.000000 496.150000 ;
        RECT 60.000000 499.850000 65.000000 500.150000 ;
        RECT 60.000000 503.850000 65.000000 504.150000 ;
        RECT 60.000000 507.850000 65.000000 508.150000 ;
        RECT 60.000000 515.850000 65.000000 516.150000 ;
        RECT 60.000000 511.850000 65.000000 512.150000 ;
        RECT 110.000000 499.850000 115.000000 500.150000 ;
        RECT 110.000000 495.850000 115.000000 496.150000 ;
        RECT 110.000000 491.850000 115.000000 492.150000 ;
        RECT 110.000000 507.850000 115.000000 508.150000 ;
        RECT 110.000000 503.850000 115.000000 504.150000 ;
        RECT 110.000000 515.850000 115.000000 516.150000 ;
        RECT 110.000000 511.850000 115.000000 512.150000 ;
        RECT 160.000000 491.850000 165.000000 492.150000 ;
        RECT 160.000000 495.850000 165.000000 496.150000 ;
        RECT 160.000000 499.850000 165.000000 500.150000 ;
        RECT 160.000000 507.850000 165.000000 508.150000 ;
        RECT 160.000000 503.850000 165.000000 504.150000 ;
        RECT 160.000000 515.850000 165.000000 516.150000 ;
        RECT 160.000000 511.850000 165.000000 512.150000 ;
        RECT 210.000000 491.850000 215.000000 492.150000 ;
        RECT 210.000000 495.850000 215.000000 496.150000 ;
        RECT 210.000000 499.850000 215.000000 500.150000 ;
        RECT 210.000000 503.850000 215.000000 504.150000 ;
        RECT 210.000000 507.850000 215.000000 508.150000 ;
        RECT 210.000000 515.850000 215.000000 516.150000 ;
        RECT 210.000000 511.850000 215.000000 512.150000 ;
        RECT 260.000000 495.850000 265.000000 496.150000 ;
        RECT 260.000000 491.850000 265.000000 492.150000 ;
        RECT 260.000000 499.850000 265.000000 500.150000 ;
        RECT 260.000000 507.850000 265.000000 508.150000 ;
        RECT 260.000000 503.850000 265.000000 504.150000 ;
        RECT 260.000000 515.850000 265.000000 516.150000 ;
        RECT 260.000000 511.850000 265.000000 512.150000 ;
        RECT 360.000000 379.850000 365.000000 380.150000 ;
        RECT 310.000000 379.850000 315.000000 380.150000 ;
        RECT 310.000000 343.850000 315.000000 344.150000 ;
        RECT 310.000000 351.850000 315.000000 352.150000 ;
        RECT 310.000000 347.850000 315.000000 348.150000 ;
        RECT 310.000000 355.850000 315.000000 356.150000 ;
        RECT 310.000000 359.850000 315.000000 360.150000 ;
        RECT 310.000000 363.850000 315.000000 364.150000 ;
        RECT 310.000000 367.850000 315.000000 368.150000 ;
        RECT 310.000000 371.850000 315.000000 372.150000 ;
        RECT 310.000000 375.850000 315.000000 376.150000 ;
        RECT 360.000000 343.850000 365.000000 344.150000 ;
        RECT 360.000000 347.850000 365.000000 348.150000 ;
        RECT 360.000000 351.850000 365.000000 352.150000 ;
        RECT 360.000000 355.850000 365.000000 356.150000 ;
        RECT 360.000000 359.850000 365.000000 360.150000 ;
        RECT 360.000000 375.850000 365.000000 376.150000 ;
        RECT 360.000000 371.850000 365.000000 372.150000 ;
        RECT 360.000000 367.850000 365.000000 368.150000 ;
        RECT 360.000000 363.850000 365.000000 364.150000 ;
        RECT 310.000000 383.850000 315.000000 384.150000 ;
        RECT 310.000000 387.850000 315.000000 388.150000 ;
        RECT 310.000000 391.850000 315.000000 392.150000 ;
        RECT 310.000000 395.850000 315.000000 396.150000 ;
        RECT 310.000000 407.850000 315.000000 408.150000 ;
        RECT 310.000000 399.850000 315.000000 400.150000 ;
        RECT 310.000000 403.850000 315.000000 404.150000 ;
        RECT 310.000000 411.850000 315.000000 412.150000 ;
        RECT 310.000000 415.850000 315.000000 416.150000 ;
        RECT 360.000000 383.850000 365.000000 384.150000 ;
        RECT 360.000000 387.850000 365.000000 388.150000 ;
        RECT 360.000000 391.850000 365.000000 392.150000 ;
        RECT 360.000000 395.850000 365.000000 396.150000 ;
        RECT 360.000000 407.850000 365.000000 408.150000 ;
        RECT 360.000000 399.850000 365.000000 400.150000 ;
        RECT 360.000000 403.850000 365.000000 404.150000 ;
        RECT 360.000000 411.850000 365.000000 412.150000 ;
        RECT 360.000000 415.850000 365.000000 416.150000 ;
        RECT 410.000000 379.850000 415.000000 380.150000 ;
        RECT 410.000000 351.850000 415.000000 352.150000 ;
        RECT 410.000000 347.850000 415.000000 348.150000 ;
        RECT 410.000000 343.850000 415.000000 344.150000 ;
        RECT 410.000000 355.850000 415.000000 356.150000 ;
        RECT 410.000000 359.850000 415.000000 360.150000 ;
        RECT 410.000000 375.850000 415.000000 376.150000 ;
        RECT 410.000000 371.850000 415.000000 372.150000 ;
        RECT 410.000000 367.850000 415.000000 368.150000 ;
        RECT 410.000000 363.850000 415.000000 364.150000 ;
        RECT 410.000000 383.850000 415.000000 384.150000 ;
        RECT 410.000000 387.850000 415.000000 388.150000 ;
        RECT 410.000000 391.850000 415.000000 392.150000 ;
        RECT 410.000000 395.850000 415.000000 396.150000 ;
        RECT 410.000000 407.850000 415.000000 408.150000 ;
        RECT 410.000000 399.850000 415.000000 400.150000 ;
        RECT 410.000000 403.850000 415.000000 404.150000 ;
        RECT 410.000000 411.850000 415.000000 412.150000 ;
        RECT 410.000000 415.850000 415.000000 416.150000 ;
        RECT 310.000000 419.850000 315.000000 420.150000 ;
        RECT 310.000000 423.850000 315.000000 424.150000 ;
        RECT 310.000000 427.850000 315.000000 428.150000 ;
        RECT 310.000000 431.850000 315.000000 432.150000 ;
        RECT 310.000000 439.850000 315.000000 440.150000 ;
        RECT 310.000000 435.850000 315.000000 436.150000 ;
        RECT 310.000000 443.850000 315.000000 444.150000 ;
        RECT 310.000000 447.850000 315.000000 448.150000 ;
        RECT 310.000000 451.850000 315.000000 452.150000 ;
        RECT 360.000000 419.850000 365.000000 420.150000 ;
        RECT 360.000000 423.850000 365.000000 424.150000 ;
        RECT 360.000000 427.850000 365.000000 428.150000 ;
        RECT 360.000000 431.850000 365.000000 432.150000 ;
        RECT 360.000000 435.850000 365.000000 436.150000 ;
        RECT 360.000000 439.850000 365.000000 440.150000 ;
        RECT 360.000000 443.850000 365.000000 444.150000 ;
        RECT 360.000000 447.850000 365.000000 448.150000 ;
        RECT 360.000000 451.850000 365.000000 452.150000 ;
        RECT 310.000000 459.850000 315.000000 460.150000 ;
        RECT 310.000000 455.850000 315.000000 456.150000 ;
        RECT 310.000000 467.850000 315.000000 468.150000 ;
        RECT 310.000000 463.850000 315.000000 464.150000 ;
        RECT 310.000000 471.850000 315.000000 472.150000 ;
        RECT 310.000000 475.850000 315.000000 476.150000 ;
        RECT 310.000000 479.850000 315.000000 480.150000 ;
        RECT 310.000000 483.850000 315.000000 484.150000 ;
        RECT 310.000000 487.850000 315.000000 488.150000 ;
        RECT 360.000000 455.850000 365.000000 456.150000 ;
        RECT 360.000000 459.850000 365.000000 460.150000 ;
        RECT 360.000000 463.850000 365.000000 464.150000 ;
        RECT 360.000000 467.850000 365.000000 468.150000 ;
        RECT 360.000000 471.850000 365.000000 472.150000 ;
        RECT 360.000000 475.850000 365.000000 476.150000 ;
        RECT 360.000000 479.850000 365.000000 480.150000 ;
        RECT 360.000000 483.850000 365.000000 484.150000 ;
        RECT 360.000000 487.850000 365.000000 488.150000 ;
        RECT 410.000000 423.850000 415.000000 424.150000 ;
        RECT 410.000000 419.850000 415.000000 420.150000 ;
        RECT 410.000000 427.850000 415.000000 428.150000 ;
        RECT 410.000000 431.850000 415.000000 432.150000 ;
        RECT 410.000000 439.850000 415.000000 440.150000 ;
        RECT 410.000000 435.850000 415.000000 436.150000 ;
        RECT 410.000000 443.850000 415.000000 444.150000 ;
        RECT 410.000000 447.850000 415.000000 448.150000 ;
        RECT 410.000000 451.850000 415.000000 452.150000 ;
        RECT 371.000000 479.850000 381.000000 480.150000 ;
        RECT 371.000000 483.850000 381.000000 484.150000 ;
        RECT 371.000000 487.850000 381.000000 488.150000 ;
        RECT 410.000000 455.850000 415.000000 456.150000 ;
        RECT 410.000000 459.850000 415.000000 460.150000 ;
        RECT 410.000000 467.850000 415.000000 468.150000 ;
        RECT 410.000000 463.850000 415.000000 464.150000 ;
        RECT 410.000000 471.850000 415.000000 472.150000 ;
        RECT 410.000000 475.850000 415.000000 476.150000 ;
        RECT 410.000000 479.850000 415.000000 480.150000 ;
        RECT 410.000000 483.850000 415.000000 484.150000 ;
        RECT 410.000000 487.850000 415.000000 488.150000 ;
        RECT 460.000000 379.850000 465.000000 380.150000 ;
        RECT 510.000000 379.850000 515.000000 380.150000 ;
        RECT 460.000000 347.850000 465.000000 348.150000 ;
        RECT 460.000000 343.850000 465.000000 344.150000 ;
        RECT 460.000000 375.850000 465.000000 376.150000 ;
        RECT 460.000000 371.850000 465.000000 372.150000 ;
        RECT 510.000000 343.850000 515.000000 344.150000 ;
        RECT 510.000000 351.850000 515.000000 352.150000 ;
        RECT 510.000000 347.850000 515.000000 348.150000 ;
        RECT 510.000000 359.850000 515.000000 360.150000 ;
        RECT 510.000000 355.850000 515.000000 356.150000 ;
        RECT 510.000000 363.850000 515.000000 364.150000 ;
        RECT 510.000000 367.850000 515.000000 368.150000 ;
        RECT 510.000000 375.850000 515.000000 376.150000 ;
        RECT 510.000000 371.850000 515.000000 372.150000 ;
        RECT 460.000000 395.850000 465.000000 396.150000 ;
        RECT 460.000000 391.850000 465.000000 392.150000 ;
        RECT 460.000000 387.850000 465.000000 388.150000 ;
        RECT 460.000000 383.850000 465.000000 384.150000 ;
        RECT 510.000000 383.850000 515.000000 384.150000 ;
        RECT 510.000000 387.850000 515.000000 388.150000 ;
        RECT 510.000000 391.850000 515.000000 392.150000 ;
        RECT 510.000000 395.850000 515.000000 396.150000 ;
        RECT 510.000000 407.850000 515.000000 408.150000 ;
        RECT 510.000000 399.850000 515.000000 400.150000 ;
        RECT 510.000000 403.850000 515.000000 404.150000 ;
        RECT 510.000000 411.850000 515.000000 412.150000 ;
        RECT 510.000000 415.850000 515.000000 416.150000 ;
        RECT 560.000000 379.850000 565.000000 380.150000 ;
        RECT 560.000000 359.850000 565.000000 360.150000 ;
        RECT 560.000000 355.850000 565.000000 356.150000 ;
        RECT 560.000000 351.850000 565.000000 352.150000 ;
        RECT 560.000000 347.850000 565.000000 348.150000 ;
        RECT 560.000000 343.850000 565.000000 344.150000 ;
        RECT 560.000000 375.850000 565.000000 376.150000 ;
        RECT 560.000000 371.850000 565.000000 372.150000 ;
        RECT 560.000000 367.850000 565.000000 368.150000 ;
        RECT 560.000000 363.850000 565.000000 364.150000 ;
        RECT 560.000000 383.850000 565.000000 384.150000 ;
        RECT 560.000000 387.850000 565.000000 388.150000 ;
        RECT 560.000000 395.850000 565.000000 396.150000 ;
        RECT 560.000000 391.850000 565.000000 392.150000 ;
        RECT 560.000000 407.850000 565.000000 408.150000 ;
        RECT 560.000000 399.850000 565.000000 400.150000 ;
        RECT 560.000000 403.850000 565.000000 404.150000 ;
        RECT 560.000000 415.850000 565.000000 416.150000 ;
        RECT 560.000000 411.850000 565.000000 412.150000 ;
        RECT 460.000000 419.850000 465.000000 420.150000 ;
        RECT 460.000000 423.850000 465.000000 424.150000 ;
        RECT 460.000000 427.850000 465.000000 428.150000 ;
        RECT 460.000000 431.850000 465.000000 432.150000 ;
        RECT 460.000000 435.850000 465.000000 436.150000 ;
        RECT 460.000000 439.850000 465.000000 440.150000 ;
        RECT 460.000000 443.850000 465.000000 444.150000 ;
        RECT 460.000000 447.850000 465.000000 448.150000 ;
        RECT 460.000000 451.850000 465.000000 452.150000 ;
        RECT 510.000000 419.850000 515.000000 420.150000 ;
        RECT 510.000000 423.850000 515.000000 424.150000 ;
        RECT 510.000000 427.850000 515.000000 428.150000 ;
        RECT 510.000000 431.850000 515.000000 432.150000 ;
        RECT 510.000000 439.850000 515.000000 440.150000 ;
        RECT 510.000000 435.850000 515.000000 436.150000 ;
        RECT 510.000000 443.850000 515.000000 444.150000 ;
        RECT 510.000000 447.850000 515.000000 448.150000 ;
        RECT 510.000000 451.850000 515.000000 452.150000 ;
        RECT 460.000000 455.850000 465.000000 456.150000 ;
        RECT 460.000000 459.850000 465.000000 460.150000 ;
        RECT 460.000000 463.850000 465.000000 464.150000 ;
        RECT 460.000000 467.850000 465.000000 468.150000 ;
        RECT 460.000000 471.850000 465.000000 472.150000 ;
        RECT 460.000000 475.850000 465.000000 476.150000 ;
        RECT 460.000000 479.850000 465.000000 480.150000 ;
        RECT 460.000000 483.850000 465.000000 484.150000 ;
        RECT 460.000000 487.850000 465.000000 488.150000 ;
        RECT 510.000000 455.850000 515.000000 456.150000 ;
        RECT 510.000000 459.850000 515.000000 460.150000 ;
        RECT 510.000000 467.850000 515.000000 468.150000 ;
        RECT 510.000000 463.850000 515.000000 464.150000 ;
        RECT 510.000000 471.850000 515.000000 472.150000 ;
        RECT 510.000000 475.850000 515.000000 476.150000 ;
        RECT 510.000000 479.850000 515.000000 480.150000 ;
        RECT 510.000000 483.850000 515.000000 484.150000 ;
        RECT 510.000000 487.850000 515.000000 488.150000 ;
        RECT 560.000000 423.850000 565.000000 424.150000 ;
        RECT 560.000000 419.850000 565.000000 420.150000 ;
        RECT 560.000000 427.850000 565.000000 428.150000 ;
        RECT 560.000000 431.850000 565.000000 432.150000 ;
        RECT 560.000000 435.850000 565.000000 436.150000 ;
        RECT 560.000000 439.850000 565.000000 440.150000 ;
        RECT 560.000000 443.850000 565.000000 444.150000 ;
        RECT 560.000000 447.850000 565.000000 448.150000 ;
        RECT 560.000000 451.850000 565.000000 452.150000 ;
        RECT 560.000000 455.850000 565.000000 456.150000 ;
        RECT 560.000000 459.850000 565.000000 460.150000 ;
        RECT 560.000000 467.850000 565.000000 468.150000 ;
        RECT 560.000000 463.850000 565.000000 464.150000 ;
        RECT 560.000000 471.850000 565.000000 472.150000 ;
        RECT 560.000000 475.850000 565.000000 476.150000 ;
        RECT 560.000000 479.850000 565.000000 480.150000 ;
        RECT 560.000000 483.850000 565.000000 484.150000 ;
        RECT 560.000000 487.850000 565.000000 488.150000 ;
        RECT 310.000000 495.850000 315.000000 496.150000 ;
        RECT 310.000000 491.850000 315.000000 492.150000 ;
        RECT 310.000000 499.850000 315.000000 500.150000 ;
        RECT 310.000000 507.850000 315.000000 508.150000 ;
        RECT 310.000000 503.850000 315.000000 504.150000 ;
        RECT 310.000000 515.850000 315.000000 516.150000 ;
        RECT 310.000000 511.850000 315.000000 512.150000 ;
        RECT 360.000000 491.850000 365.000000 492.150000 ;
        RECT 360.000000 495.850000 365.000000 496.150000 ;
        RECT 360.000000 499.850000 365.000000 500.150000 ;
        RECT 360.000000 503.850000 365.000000 504.150000 ;
        RECT 360.000000 507.850000 365.000000 508.150000 ;
        RECT 360.000000 511.850000 365.000000 512.150000 ;
        RECT 360.000000 515.850000 365.000000 516.150000 ;
        RECT 360.000000 519.850000 365.000000 520.150000 ;
        RECT 360.000000 523.850000 365.000000 524.150000 ;
        RECT 360.000000 527.850000 365.000000 528.150000 ;
        RECT 360.000000 531.850000 365.000000 532.150000 ;
        RECT 360.000000 535.850000 365.000000 536.150000 ;
        RECT 360.000000 539.850000 365.000000 540.150000 ;
        RECT 360.000000 543.850000 365.000000 544.150000 ;
        RECT 360.000000 555.850000 365.000000 556.150000 ;
        RECT 360.000000 547.850000 365.000000 548.150000 ;
        RECT 360.000000 551.850000 365.000000 552.150000 ;
        RECT 360.000000 559.850000 365.000000 560.150000 ;
        RECT 360.000000 563.850000 365.000000 564.150000 ;
        RECT 371.000000 491.850000 381.000000 492.150000 ;
        RECT 371.000000 495.850000 381.000000 496.150000 ;
        RECT 371.000000 499.850000 381.000000 500.150000 ;
        RECT 371.000000 503.850000 381.000000 504.150000 ;
        RECT 371.000000 507.850000 381.000000 508.150000 ;
        RECT 371.000000 511.850000 381.000000 512.150000 ;
        RECT 371.000000 515.850000 381.000000 516.150000 ;
        RECT 371.000000 519.850000 381.000000 520.150000 ;
        RECT 371.000000 523.850000 381.000000 524.150000 ;
        RECT 371.000000 527.850000 381.000000 528.150000 ;
        RECT 410.000000 495.850000 415.000000 496.150000 ;
        RECT 410.000000 491.850000 415.000000 492.150000 ;
        RECT 410.000000 499.850000 415.000000 500.150000 ;
        RECT 410.000000 503.850000 415.000000 504.150000 ;
        RECT 371.000000 531.850000 381.000000 532.150000 ;
        RECT 371.000000 535.850000 381.000000 536.150000 ;
        RECT 371.000000 539.850000 381.000000 540.150000 ;
        RECT 371.000000 543.850000 381.000000 544.150000 ;
        RECT 371.000000 555.850000 381.000000 556.150000 ;
        RECT 371.000000 547.850000 381.000000 548.150000 ;
        RECT 371.000000 551.850000 381.000000 552.150000 ;
        RECT 371.000000 559.850000 381.000000 560.150000 ;
        RECT 371.000000 563.850000 381.000000 564.150000 ;
        RECT 360.000000 583.850000 365.000000 584.150000 ;
        RECT 360.000000 567.850000 365.000000 568.150000 ;
        RECT 360.000000 571.850000 365.000000 572.150000 ;
        RECT 360.000000 575.850000 365.000000 576.150000 ;
        RECT 360.000000 579.850000 365.000000 580.150000 ;
        RECT 360.000000 587.850000 365.000000 588.150000 ;
        RECT 360.000000 591.850000 365.000000 592.150000 ;
        RECT 360.000000 595.850000 365.000000 596.150000 ;
        RECT 360.000000 599.850000 365.000000 600.150000 ;
        RECT 360.000000 603.850000 365.000000 604.150000 ;
        RECT 360.000000 607.850000 365.000000 608.150000 ;
        RECT 360.000000 611.850000 365.000000 612.150000 ;
        RECT 360.000000 615.850000 365.000000 616.150000 ;
        RECT 360.000000 619.850000 365.000000 620.150000 ;
        RECT 360.000000 623.850000 365.000000 624.150000 ;
        RECT 360.000000 627.850000 365.000000 628.150000 ;
        RECT 360.000000 631.850000 365.000000 632.150000 ;
        RECT 360.000000 635.850000 365.000000 636.150000 ;
        RECT 371.000000 583.850000 381.000000 584.150000 ;
        RECT 371.000000 579.850000 381.000000 580.150000 ;
        RECT 371.000000 575.850000 381.000000 576.150000 ;
        RECT 371.000000 571.850000 381.000000 572.150000 ;
        RECT 371.000000 567.850000 381.000000 568.150000 ;
        RECT 371.000000 587.850000 381.000000 588.150000 ;
        RECT 371.000000 591.850000 381.000000 592.150000 ;
        RECT 371.000000 595.850000 381.000000 596.150000 ;
        RECT 371.000000 599.850000 381.000000 600.150000 ;
        RECT 371.000000 603.850000 381.000000 604.150000 ;
        RECT 371.000000 607.850000 381.000000 608.150000 ;
        RECT 371.000000 611.850000 381.000000 612.150000 ;
        RECT 371.000000 615.850000 381.000000 616.150000 ;
        RECT 371.000000 619.850000 381.000000 620.150000 ;
        RECT 371.000000 635.850000 381.000000 636.150000 ;
        RECT 371.000000 631.850000 381.000000 632.150000 ;
        RECT 371.000000 627.850000 381.000000 628.150000 ;
        RECT 371.000000 623.850000 381.000000 624.150000 ;
        RECT 460.000000 495.850000 465.000000 496.150000 ;
        RECT 460.000000 491.850000 465.000000 492.150000 ;
        RECT 460.000000 499.850000 465.000000 500.150000 ;
        RECT 460.000000 503.850000 465.000000 504.150000 ;
        RECT 510.000000 495.850000 515.000000 496.150000 ;
        RECT 510.000000 491.850000 515.000000 492.150000 ;
        RECT 510.000000 499.850000 515.000000 500.150000 ;
        RECT 510.000000 503.850000 515.000000 504.150000 ;
        RECT 560.000000 503.850000 565.000000 504.150000 ;
        RECT 560.000000 499.850000 565.000000 500.150000 ;
        RECT 560.000000 495.850000 565.000000 496.150000 ;
        RECT 560.000000 491.850000 565.000000 492.150000 ;
        RECT 360.000000 639.850000 365.000000 640.150000 ;
        RECT 360.000000 643.850000 365.000000 644.150000 ;
        RECT 360.000000 647.850000 365.000000 648.150000 ;
        RECT 360.000000 651.850000 365.000000 652.150000 ;
        RECT 360.000000 655.850000 365.000000 656.150000 ;
        RECT 360.000000 659.850000 365.000000 660.150000 ;
        RECT 360.000000 663.850000 365.000000 664.150000 ;
        RECT 360.000000 667.850000 365.000000 668.150000 ;
        RECT 360.000000 671.850000 365.000000 672.150000 ;
        RECT 360.000000 675.850000 365.000000 676.150000 ;
        RECT 310.000000 679.850000 315.000000 680.150000 ;
        RECT 310.000000 683.850000 315.000000 684.150000 ;
        RECT 360.000000 679.850000 365.000000 680.150000 ;
        RECT 360.000000 683.850000 365.000000 684.150000 ;
        RECT 371.000000 639.850000 381.000000 640.150000 ;
        RECT 371.000000 643.850000 381.000000 644.150000 ;
        RECT 371.000000 647.850000 381.000000 648.150000 ;
        RECT 371.000000 651.850000 381.000000 652.150000 ;
        RECT 371.000000 655.850000 381.000000 656.150000 ;
        RECT 371.000000 667.850000 381.000000 668.150000 ;
        RECT 371.000000 663.850000 381.000000 664.150000 ;
        RECT 371.000000 659.850000 381.000000 660.150000 ;
        RECT 410.000000 659.850000 415.000000 660.150000 ;
        RECT 410.000000 663.850000 415.000000 664.150000 ;
        RECT 410.000000 667.850000 415.000000 668.150000 ;
        RECT 410.000000 671.850000 415.000000 672.150000 ;
        RECT 410.000000 675.850000 415.000000 676.150000 ;
        RECT 410.000000 683.850000 415.000000 684.150000 ;
        RECT 410.000000 679.850000 415.000000 680.150000 ;
        RECT 460.000000 659.850000 465.000000 660.150000 ;
        RECT 460.000000 663.850000 465.000000 664.150000 ;
        RECT 460.000000 667.850000 465.000000 668.150000 ;
        RECT 460.000000 671.850000 465.000000 672.150000 ;
        RECT 460.000000 675.850000 465.000000 676.150000 ;
        RECT 510.000000 659.850000 515.000000 660.150000 ;
        RECT 510.000000 663.850000 515.000000 664.150000 ;
        RECT 510.000000 667.850000 515.000000 668.150000 ;
        RECT 510.000000 671.850000 515.000000 672.150000 ;
        RECT 510.000000 675.850000 515.000000 676.150000 ;
        RECT 460.000000 683.850000 465.000000 684.150000 ;
        RECT 460.000000 679.850000 465.000000 680.150000 ;
        RECT 510.000000 683.850000 515.000000 684.150000 ;
        RECT 510.000000 679.850000 515.000000 680.150000 ;
        RECT 560.000000 659.850000 565.000000 660.150000 ;
        RECT 560.000000 663.850000 565.000000 664.150000 ;
        RECT 560.000000 667.850000 565.000000 668.150000 ;
        RECT 560.000000 671.850000 565.000000 672.150000 ;
        RECT 560.000000 675.850000 565.000000 676.150000 ;
        RECT 560.000000 683.850000 565.000000 684.150000 ;
        RECT 560.000000 679.850000 565.000000 680.150000 ;
        RECT 610.000000 379.850000 615.000000 380.150000 ;
        RECT 660.000000 379.850000 665.000000 380.150000 ;
        RECT 610.000000 343.850000 615.000000 344.150000 ;
        RECT 610.000000 347.850000 615.000000 348.150000 ;
        RECT 610.000000 351.850000 615.000000 352.150000 ;
        RECT 610.000000 355.850000 615.000000 356.150000 ;
        RECT 610.000000 359.850000 615.000000 360.150000 ;
        RECT 610.000000 375.850000 615.000000 376.150000 ;
        RECT 610.000000 371.850000 615.000000 372.150000 ;
        RECT 610.000000 367.850000 615.000000 368.150000 ;
        RECT 610.000000 363.850000 615.000000 364.150000 ;
        RECT 660.000000 343.850000 665.000000 344.150000 ;
        RECT 660.000000 347.850000 665.000000 348.150000 ;
        RECT 660.000000 351.850000 665.000000 352.150000 ;
        RECT 660.000000 359.850000 665.000000 360.150000 ;
        RECT 660.000000 355.850000 665.000000 356.150000 ;
        RECT 660.000000 363.850000 665.000000 364.150000 ;
        RECT 660.000000 367.850000 665.000000 368.150000 ;
        RECT 660.000000 371.850000 665.000000 372.150000 ;
        RECT 660.000000 375.850000 665.000000 376.150000 ;
        RECT 610.000000 383.850000 615.000000 384.150000 ;
        RECT 610.000000 387.850000 615.000000 388.150000 ;
        RECT 610.000000 391.850000 615.000000 392.150000 ;
        RECT 610.000000 395.850000 615.000000 396.150000 ;
        RECT 610.000000 407.850000 615.000000 408.150000 ;
        RECT 610.000000 399.850000 615.000000 400.150000 ;
        RECT 610.000000 403.850000 615.000000 404.150000 ;
        RECT 610.000000 411.850000 615.000000 412.150000 ;
        RECT 610.000000 415.850000 615.000000 416.150000 ;
        RECT 660.000000 383.850000 665.000000 384.150000 ;
        RECT 660.000000 387.850000 665.000000 388.150000 ;
        RECT 660.000000 391.850000 665.000000 392.150000 ;
        RECT 660.000000 395.850000 665.000000 396.150000 ;
        RECT 660.000000 407.850000 665.000000 408.150000 ;
        RECT 660.000000 399.850000 665.000000 400.150000 ;
        RECT 660.000000 403.850000 665.000000 404.150000 ;
        RECT 660.000000 411.850000 665.000000 412.150000 ;
        RECT 660.000000 415.850000 665.000000 416.150000 ;
        RECT 710.000000 379.850000 715.000000 380.150000 ;
        RECT 710.000000 359.850000 715.000000 360.150000 ;
        RECT 710.000000 355.850000 715.000000 356.150000 ;
        RECT 710.000000 351.850000 715.000000 352.150000 ;
        RECT 710.000000 347.850000 715.000000 348.150000 ;
        RECT 710.000000 343.850000 715.000000 344.150000 ;
        RECT 710.000000 375.850000 715.000000 376.150000 ;
        RECT 710.000000 371.850000 715.000000 372.150000 ;
        RECT 710.000000 367.850000 715.000000 368.150000 ;
        RECT 710.000000 363.850000 715.000000 364.150000 ;
        RECT 710.000000 383.850000 715.000000 384.150000 ;
        RECT 710.000000 387.850000 715.000000 388.150000 ;
        RECT 710.000000 391.850000 715.000000 392.150000 ;
        RECT 710.000000 395.850000 715.000000 396.150000 ;
        RECT 710.000000 407.850000 715.000000 408.150000 ;
        RECT 710.000000 403.850000 715.000000 404.150000 ;
        RECT 710.000000 399.850000 715.000000 400.150000 ;
        RECT 710.000000 415.850000 715.000000 416.150000 ;
        RECT 710.000000 411.850000 715.000000 412.150000 ;
        RECT 610.000000 419.850000 615.000000 420.150000 ;
        RECT 610.000000 423.850000 615.000000 424.150000 ;
        RECT 610.000000 427.850000 615.000000 428.150000 ;
        RECT 610.000000 431.850000 615.000000 432.150000 ;
        RECT 610.000000 435.850000 615.000000 436.150000 ;
        RECT 610.000000 439.850000 615.000000 440.150000 ;
        RECT 610.000000 443.850000 615.000000 444.150000 ;
        RECT 610.000000 447.850000 615.000000 448.150000 ;
        RECT 610.000000 451.850000 615.000000 452.150000 ;
        RECT 660.000000 419.850000 665.000000 420.150000 ;
        RECT 660.000000 423.850000 665.000000 424.150000 ;
        RECT 660.000000 427.850000 665.000000 428.150000 ;
        RECT 660.000000 431.850000 665.000000 432.150000 ;
        RECT 660.000000 435.850000 665.000000 436.150000 ;
        RECT 660.000000 439.850000 665.000000 440.150000 ;
        RECT 660.000000 443.850000 665.000000 444.150000 ;
        RECT 660.000000 447.850000 665.000000 448.150000 ;
        RECT 660.000000 451.850000 665.000000 452.150000 ;
        RECT 610.000000 455.850000 615.000000 456.150000 ;
        RECT 610.000000 459.850000 615.000000 460.150000 ;
        RECT 610.000000 463.850000 615.000000 464.150000 ;
        RECT 610.000000 467.850000 615.000000 468.150000 ;
        RECT 610.000000 471.850000 615.000000 472.150000 ;
        RECT 610.000000 487.850000 615.000000 488.150000 ;
        RECT 610.000000 483.850000 615.000000 484.150000 ;
        RECT 610.000000 479.850000 615.000000 480.150000 ;
        RECT 610.000000 475.850000 615.000000 476.150000 ;
        RECT 660.000000 455.850000 665.000000 456.150000 ;
        RECT 660.000000 459.850000 665.000000 460.150000 ;
        RECT 660.000000 463.850000 665.000000 464.150000 ;
        RECT 660.000000 467.850000 665.000000 468.150000 ;
        RECT 660.000000 471.850000 665.000000 472.150000 ;
        RECT 660.000000 479.850000 665.000000 480.150000 ;
        RECT 660.000000 475.850000 665.000000 476.150000 ;
        RECT 660.000000 487.850000 665.000000 488.150000 ;
        RECT 660.000000 483.850000 665.000000 484.150000 ;
        RECT 721.000000 431.850000 731.000000 432.150000 ;
        RECT 721.000000 419.850000 731.000000 420.150000 ;
        RECT 721.000000 423.850000 731.000000 424.150000 ;
        RECT 721.000000 427.850000 731.000000 428.150000 ;
        RECT 710.000000 419.850000 715.000000 420.150000 ;
        RECT 710.000000 423.850000 715.000000 424.150000 ;
        RECT 710.000000 427.850000 715.000000 428.150000 ;
        RECT 710.000000 431.850000 715.000000 432.150000 ;
        RECT 721.000000 435.850000 731.000000 436.150000 ;
        RECT 721.000000 439.850000 731.000000 440.150000 ;
        RECT 721.000000 443.850000 731.000000 444.150000 ;
        RECT 721.000000 447.850000 731.000000 448.150000 ;
        RECT 721.000000 451.850000 731.000000 452.150000 ;
        RECT 710.000000 439.850000 715.000000 440.150000 ;
        RECT 710.000000 435.850000 715.000000 436.150000 ;
        RECT 710.000000 443.850000 715.000000 444.150000 ;
        RECT 710.000000 447.850000 715.000000 448.150000 ;
        RECT 710.000000 451.850000 715.000000 452.150000 ;
        RECT 721.000000 459.850000 731.000000 460.150000 ;
        RECT 721.000000 455.850000 731.000000 456.150000 ;
        RECT 721.000000 463.850000 731.000000 464.150000 ;
        RECT 721.000000 467.850000 731.000000 468.150000 ;
        RECT 721.000000 471.850000 731.000000 472.150000 ;
        RECT 710.000000 455.850000 715.000000 456.150000 ;
        RECT 710.000000 459.850000 715.000000 460.150000 ;
        RECT 710.000000 463.850000 715.000000 464.150000 ;
        RECT 710.000000 467.850000 715.000000 468.150000 ;
        RECT 710.000000 471.850000 715.000000 472.150000 ;
        RECT 721.000000 487.850000 731.000000 488.150000 ;
        RECT 721.000000 483.850000 731.000000 484.150000 ;
        RECT 721.000000 479.850000 731.000000 480.150000 ;
        RECT 721.000000 475.850000 731.000000 476.150000 ;
        RECT 710.000000 487.850000 715.000000 488.150000 ;
        RECT 710.000000 483.850000 715.000000 484.150000 ;
        RECT 710.000000 475.850000 715.000000 476.150000 ;
        RECT 710.000000 479.850000 715.000000 480.150000 ;
        RECT 810.000000 379.850000 815.000000 380.150000 ;
        RECT 760.000000 379.850000 765.000000 380.150000 ;
        RECT 760.000000 343.850000 765.000000 344.150000 ;
        RECT 760.000000 347.850000 765.000000 348.150000 ;
        RECT 760.000000 351.850000 765.000000 352.150000 ;
        RECT 760.000000 355.850000 765.000000 356.150000 ;
        RECT 760.000000 359.850000 765.000000 360.150000 ;
        RECT 760.000000 375.850000 765.000000 376.150000 ;
        RECT 760.000000 371.850000 765.000000 372.150000 ;
        RECT 760.000000 367.850000 765.000000 368.150000 ;
        RECT 760.000000 363.850000 765.000000 364.150000 ;
        RECT 810.000000 343.850000 815.000000 344.150000 ;
        RECT 810.000000 347.850000 815.000000 348.150000 ;
        RECT 810.000000 351.850000 815.000000 352.150000 ;
        RECT 810.000000 359.850000 815.000000 360.150000 ;
        RECT 810.000000 355.850000 815.000000 356.150000 ;
        RECT 810.000000 363.850000 815.000000 364.150000 ;
        RECT 810.000000 367.850000 815.000000 368.150000 ;
        RECT 810.000000 375.850000 815.000000 376.150000 ;
        RECT 810.000000 371.850000 815.000000 372.150000 ;
        RECT 760.000000 383.850000 765.000000 384.150000 ;
        RECT 760.000000 387.850000 765.000000 388.150000 ;
        RECT 760.000000 391.850000 765.000000 392.150000 ;
        RECT 760.000000 395.850000 765.000000 396.150000 ;
        RECT 760.000000 407.850000 765.000000 408.150000 ;
        RECT 760.000000 399.850000 765.000000 400.150000 ;
        RECT 760.000000 403.850000 765.000000 404.150000 ;
        RECT 760.000000 411.850000 765.000000 412.150000 ;
        RECT 760.000000 415.850000 765.000000 416.150000 ;
        RECT 810.000000 387.850000 815.000000 388.150000 ;
        RECT 810.000000 383.850000 815.000000 384.150000 ;
        RECT 810.000000 391.850000 815.000000 392.150000 ;
        RECT 810.000000 395.850000 815.000000 396.150000 ;
        RECT 810.000000 407.850000 815.000000 408.150000 ;
        RECT 810.000000 399.850000 815.000000 400.150000 ;
        RECT 810.000000 403.850000 815.000000 404.150000 ;
        RECT 810.000000 415.850000 815.000000 416.150000 ;
        RECT 810.000000 411.850000 815.000000 412.150000 ;
        RECT 860.000000 379.850000 865.000000 380.150000 ;
        RECT 860.000000 359.850000 865.000000 360.150000 ;
        RECT 860.000000 355.850000 865.000000 356.150000 ;
        RECT 860.000000 351.850000 865.000000 352.150000 ;
        RECT 860.000000 347.850000 865.000000 348.150000 ;
        RECT 860.000000 343.850000 865.000000 344.150000 ;
        RECT 860.000000 375.850000 865.000000 376.150000 ;
        RECT 860.000000 371.850000 865.000000 372.150000 ;
        RECT 860.000000 367.850000 865.000000 368.150000 ;
        RECT 860.000000 363.850000 865.000000 364.150000 ;
        RECT 860.000000 383.850000 865.000000 384.150000 ;
        RECT 860.000000 387.850000 865.000000 388.150000 ;
        RECT 860.000000 391.850000 865.000000 392.150000 ;
        RECT 860.000000 395.850000 865.000000 396.150000 ;
        RECT 860.000000 407.850000 865.000000 408.150000 ;
        RECT 860.000000 403.850000 865.000000 404.150000 ;
        RECT 860.000000 399.850000 865.000000 400.150000 ;
        RECT 860.000000 415.850000 865.000000 416.150000 ;
        RECT 860.000000 411.850000 865.000000 412.150000 ;
        RECT 760.000000 419.850000 765.000000 420.150000 ;
        RECT 760.000000 423.850000 765.000000 424.150000 ;
        RECT 760.000000 427.850000 765.000000 428.150000 ;
        RECT 760.000000 431.850000 765.000000 432.150000 ;
        RECT 760.000000 435.850000 765.000000 436.150000 ;
        RECT 760.000000 439.850000 765.000000 440.150000 ;
        RECT 760.000000 443.850000 765.000000 444.150000 ;
        RECT 810.000000 419.850000 815.000000 420.150000 ;
        RECT 810.000000 423.850000 815.000000 424.150000 ;
        RECT 810.000000 427.850000 815.000000 428.150000 ;
        RECT 810.000000 431.850000 815.000000 432.150000 ;
        RECT 810.000000 435.850000 815.000000 436.150000 ;
        RECT 810.000000 439.850000 815.000000 440.150000 ;
        RECT 810.000000 443.850000 815.000000 444.150000 ;
        RECT 860.000000 419.850000 865.000000 420.150000 ;
        RECT 860.000000 423.850000 865.000000 424.150000 ;
        RECT 860.000000 427.850000 865.000000 428.150000 ;
        RECT 860.000000 431.850000 865.000000 432.150000 ;
        RECT 860.000000 443.850000 865.000000 444.150000 ;
        RECT 860.000000 439.850000 865.000000 440.150000 ;
        RECT 860.000000 435.850000 865.000000 436.150000 ;
        RECT 610.000000 503.850000 615.000000 504.150000 ;
        RECT 610.000000 499.850000 615.000000 500.150000 ;
        RECT 610.000000 491.850000 615.000000 492.150000 ;
        RECT 610.000000 495.850000 615.000000 496.150000 ;
        RECT 660.000000 495.850000 665.000000 496.150000 ;
        RECT 660.000000 491.850000 665.000000 492.150000 ;
        RECT 660.000000 499.850000 665.000000 500.150000 ;
        RECT 660.000000 503.850000 665.000000 504.150000 ;
        RECT 710.000000 503.850000 715.000000 504.150000 ;
        RECT 710.000000 499.850000 715.000000 500.150000 ;
        RECT 710.000000 495.850000 715.000000 496.150000 ;
        RECT 710.000000 491.850000 715.000000 492.150000 ;
        RECT 960.000000 379.850000 965.000000 380.150000 ;
        RECT 960.000000 343.850000 965.000000 344.150000 ;
        RECT 960.000000 347.850000 965.000000 348.150000 ;
        RECT 960.000000 351.850000 965.000000 352.150000 ;
        RECT 960.000000 359.850000 965.000000 360.150000 ;
        RECT 960.000000 355.850000 965.000000 356.150000 ;
        RECT 960.000000 375.850000 965.000000 376.150000 ;
        RECT 960.000000 371.850000 965.000000 372.150000 ;
        RECT 960.000000 367.850000 965.000000 368.150000 ;
        RECT 960.000000 363.850000 965.000000 364.150000 ;
        RECT 960.000000 383.850000 965.000000 384.150000 ;
        RECT 960.000000 387.850000 965.000000 388.150000 ;
        RECT 960.000000 391.850000 965.000000 392.150000 ;
        RECT 960.000000 395.850000 965.000000 396.150000 ;
        RECT 960.000000 407.850000 965.000000 408.150000 ;
        RECT 960.000000 399.850000 965.000000 400.150000 ;
        RECT 960.000000 403.850000 965.000000 404.150000 ;
        RECT 960.000000 411.850000 965.000000 412.150000 ;
        RECT 960.000000 415.850000 965.000000 416.150000 ;
        RECT 910.000000 379.850000 915.000000 380.150000 ;
        RECT 910.000000 343.850000 915.000000 344.150000 ;
        RECT 910.000000 347.850000 915.000000 348.150000 ;
        RECT 910.000000 351.850000 915.000000 352.150000 ;
        RECT 910.000000 355.850000 915.000000 356.150000 ;
        RECT 910.000000 359.850000 915.000000 360.150000 ;
        RECT 910.000000 375.850000 915.000000 376.150000 ;
        RECT 910.000000 371.850000 915.000000 372.150000 ;
        RECT 910.000000 367.850000 915.000000 368.150000 ;
        RECT 910.000000 363.850000 915.000000 364.150000 ;
        RECT 910.000000 383.850000 915.000000 384.150000 ;
        RECT 910.000000 387.850000 915.000000 388.150000 ;
        RECT 910.000000 391.850000 915.000000 392.150000 ;
        RECT 910.000000 395.850000 915.000000 396.150000 ;
        RECT 910.000000 407.850000 915.000000 408.150000 ;
        RECT 910.000000 399.850000 915.000000 400.150000 ;
        RECT 910.000000 403.850000 915.000000 404.150000 ;
        RECT 910.000000 411.850000 915.000000 412.150000 ;
        RECT 910.000000 415.850000 915.000000 416.150000 ;
        RECT 1010.000000 379.850000 1015.000000 380.150000 ;
        RECT 1010.000000 343.850000 1015.000000 344.150000 ;
        RECT 1010.000000 347.850000 1015.000000 348.150000 ;
        RECT 1010.000000 351.850000 1015.000000 352.150000 ;
        RECT 1010.000000 359.850000 1015.000000 360.150000 ;
        RECT 1010.000000 355.850000 1015.000000 356.150000 ;
        RECT 1010.000000 363.850000 1015.000000 364.150000 ;
        RECT 1010.000000 367.850000 1015.000000 368.150000 ;
        RECT 1010.000000 375.850000 1015.000000 376.150000 ;
        RECT 1010.000000 371.850000 1015.000000 372.150000 ;
        RECT 1010.000000 387.850000 1015.000000 388.150000 ;
        RECT 1010.000000 383.850000 1015.000000 384.150000 ;
        RECT 1010.000000 391.850000 1015.000000 392.150000 ;
        RECT 1010.000000 395.850000 1015.000000 396.150000 ;
        RECT 1010.000000 407.850000 1015.000000 408.150000 ;
        RECT 1010.000000 403.850000 1015.000000 404.150000 ;
        RECT 1010.000000 399.850000 1015.000000 400.150000 ;
        RECT 1010.000000 415.850000 1015.000000 416.150000 ;
        RECT 1010.000000 411.850000 1015.000000 412.150000 ;
        RECT 960.000000 431.850000 965.000000 432.150000 ;
        RECT 960.000000 427.850000 965.000000 428.150000 ;
        RECT 960.000000 423.850000 965.000000 424.150000 ;
        RECT 960.000000 419.850000 965.000000 420.150000 ;
        RECT 960.000000 443.850000 965.000000 444.150000 ;
        RECT 960.000000 439.850000 965.000000 440.150000 ;
        RECT 960.000000 435.850000 965.000000 436.150000 ;
        RECT 910.000000 419.850000 915.000000 420.150000 ;
        RECT 910.000000 423.850000 915.000000 424.150000 ;
        RECT 910.000000 427.850000 915.000000 428.150000 ;
        RECT 910.000000 431.850000 915.000000 432.150000 ;
        RECT 910.000000 435.850000 915.000000 436.150000 ;
        RECT 910.000000 439.850000 915.000000 440.150000 ;
        RECT 910.000000 443.850000 915.000000 444.150000 ;
        RECT 1010.000000 419.850000 1015.000000 420.150000 ;
        RECT 1010.000000 423.850000 1015.000000 424.150000 ;
        RECT 1010.000000 427.850000 1015.000000 428.150000 ;
        RECT 1010.000000 431.850000 1015.000000 432.150000 ;
        RECT 1010.000000 439.850000 1015.000000 440.150000 ;
        RECT 1010.000000 435.850000 1015.000000 436.150000 ;
        RECT 1010.000000 443.850000 1015.000000 444.150000 ;
        RECT 1110.000000 379.850000 1115.000000 380.150000 ;
        RECT 1110.000000 343.850000 1115.000000 344.150000 ;
        RECT 1110.000000 347.850000 1115.000000 348.150000 ;
        RECT 1110.000000 351.850000 1115.000000 352.150000 ;
        RECT 1110.000000 359.850000 1115.000000 360.150000 ;
        RECT 1110.000000 355.850000 1115.000000 356.150000 ;
        RECT 1110.000000 375.850000 1115.000000 376.150000 ;
        RECT 1110.000000 371.850000 1115.000000 372.150000 ;
        RECT 1110.000000 367.850000 1115.000000 368.150000 ;
        RECT 1110.000000 363.850000 1115.000000 364.150000 ;
        RECT 1110.000000 383.850000 1115.000000 384.150000 ;
        RECT 1110.000000 387.850000 1115.000000 388.150000 ;
        RECT 1110.000000 391.850000 1115.000000 392.150000 ;
        RECT 1110.000000 395.850000 1115.000000 396.150000 ;
        RECT 1110.000000 407.850000 1115.000000 408.150000 ;
        RECT 1110.000000 399.850000 1115.000000 400.150000 ;
        RECT 1110.000000 403.850000 1115.000000 404.150000 ;
        RECT 1110.000000 411.850000 1115.000000 412.150000 ;
        RECT 1110.000000 415.850000 1115.000000 416.150000 ;
        RECT 1060.000000 379.850000 1065.000000 380.150000 ;
        RECT 1060.000000 343.850000 1065.000000 344.150000 ;
        RECT 1060.000000 347.850000 1065.000000 348.150000 ;
        RECT 1060.000000 351.850000 1065.000000 352.150000 ;
        RECT 1060.000000 355.850000 1065.000000 356.150000 ;
        RECT 1060.000000 359.850000 1065.000000 360.150000 ;
        RECT 1060.000000 375.850000 1065.000000 376.150000 ;
        RECT 1060.000000 371.850000 1065.000000 372.150000 ;
        RECT 1060.000000 367.850000 1065.000000 368.150000 ;
        RECT 1060.000000 363.850000 1065.000000 364.150000 ;
        RECT 1060.000000 395.850000 1065.000000 396.150000 ;
        RECT 1060.000000 391.850000 1065.000000 392.150000 ;
        RECT 1060.000000 387.850000 1065.000000 388.150000 ;
        RECT 1060.000000 383.850000 1065.000000 384.150000 ;
        RECT 1060.000000 407.850000 1065.000000 408.150000 ;
        RECT 1060.000000 403.850000 1065.000000 404.150000 ;
        RECT 1060.000000 399.850000 1065.000000 400.150000 ;
        RECT 1060.000000 411.850000 1065.000000 412.150000 ;
        RECT 1060.000000 415.850000 1065.000000 416.150000 ;
        RECT 1158.000000 379.850000 1168.000000 380.150000 ;
        RECT 1158.000000 343.850000 1168.000000 344.150000 ;
        RECT 1158.000000 347.850000 1168.000000 348.150000 ;
        RECT 1158.000000 351.850000 1168.000000 352.150000 ;
        RECT 1158.000000 355.850000 1168.000000 356.150000 ;
        RECT 1158.000000 359.850000 1168.000000 360.150000 ;
        RECT 1158.000000 375.850000 1168.000000 376.150000 ;
        RECT 1158.000000 371.850000 1168.000000 372.150000 ;
        RECT 1158.000000 367.850000 1168.000000 368.150000 ;
        RECT 1158.000000 363.850000 1168.000000 364.150000 ;
        RECT 1158.000000 395.850000 1168.000000 396.150000 ;
        RECT 1158.000000 391.850000 1168.000000 392.150000 ;
        RECT 1158.000000 387.850000 1168.000000 388.150000 ;
        RECT 1158.000000 383.850000 1168.000000 384.150000 ;
        RECT 1158.000000 407.850000 1168.000000 408.150000 ;
        RECT 1158.000000 399.850000 1168.000000 400.150000 ;
        RECT 1158.000000 403.850000 1168.000000 404.150000 ;
        RECT 1158.000000 411.850000 1168.000000 412.150000 ;
        RECT 1158.000000 415.850000 1168.000000 416.150000 ;
        RECT 1110.000000 431.850000 1115.000000 432.150000 ;
        RECT 1110.000000 427.850000 1115.000000 428.150000 ;
        RECT 1110.000000 423.850000 1115.000000 424.150000 ;
        RECT 1110.000000 419.850000 1115.000000 420.150000 ;
        RECT 1110.000000 443.850000 1115.000000 444.150000 ;
        RECT 1110.000000 439.850000 1115.000000 440.150000 ;
        RECT 1110.000000 435.850000 1115.000000 436.150000 ;
        RECT 1060.000000 419.850000 1065.000000 420.150000 ;
        RECT 1060.000000 423.850000 1065.000000 424.150000 ;
        RECT 1060.000000 431.850000 1065.000000 432.150000 ;
        RECT 1060.000000 427.850000 1065.000000 428.150000 ;
        RECT 1060.000000 435.850000 1065.000000 436.150000 ;
        RECT 1060.000000 439.850000 1065.000000 440.150000 ;
        RECT 1060.000000 443.850000 1065.000000 444.150000 ;
        RECT 1158.000000 427.850000 1168.000000 428.150000 ;
        RECT 1158.000000 423.850000 1168.000000 424.150000 ;
        RECT 1158.000000 419.850000 1168.000000 420.150000 ;
        RECT 1160.000000 431.850000 1165.000000 432.150000 ;
        RECT 1160.000000 435.850000 1165.000000 436.150000 ;
        RECT 1160.000000 439.850000 1165.000000 440.150000 ;
        RECT 1160.000000 443.850000 1165.000000 444.150000 ;
        RECT 1160.000000 447.850000 1165.000000 448.150000 ;
        RECT 1160.000000 451.850000 1165.000000 452.150000 ;
        RECT 1160.000000 459.850000 1165.000000 460.150000 ;
        RECT 1160.000000 455.850000 1165.000000 456.150000 ;
        RECT 1160.000000 463.850000 1165.000000 464.150000 ;
        RECT 1160.000000 467.850000 1165.000000 468.150000 ;
        RECT 1160.000000 471.850000 1165.000000 472.150000 ;
        RECT 1160.000000 479.850000 1165.000000 480.150000 ;
        RECT 1160.000000 475.850000 1165.000000 476.150000 ;
        RECT 1160.000000 487.850000 1165.000000 488.150000 ;
        RECT 1160.000000 483.850000 1165.000000 484.150000 ;
        RECT 1160.000000 491.850000 1165.000000 492.150000 ;
        RECT 1160.000000 495.850000 1165.000000 496.150000 ;
        RECT 1160.000000 499.850000 1165.000000 500.150000 ;
        RECT 1160.000000 507.850000 1165.000000 508.150000 ;
        RECT 1160.000000 503.850000 1165.000000 504.150000 ;
        RECT 1160.000000 511.850000 1165.000000 512.150000 ;
        RECT 1160.000000 515.850000 1165.000000 516.150000 ;
        RECT 1160.000000 519.850000 1165.000000 520.150000 ;
        RECT 1160.000000 523.850000 1165.000000 524.150000 ;
        RECT 1160.000000 527.850000 1165.000000 528.150000 ;
        RECT 1160.000000 535.850000 1165.000000 536.150000 ;
        RECT 1160.000000 531.850000 1165.000000 532.150000 ;
        RECT 1160.000000 539.850000 1165.000000 540.150000 ;
        RECT 1160.000000 543.850000 1165.000000 544.150000 ;
        RECT 1160.000000 555.850000 1165.000000 556.150000 ;
        RECT 1160.000000 551.850000 1165.000000 552.150000 ;
        RECT 1160.000000 547.850000 1165.000000 548.150000 ;
        RECT 1160.000000 563.850000 1165.000000 564.150000 ;
        RECT 1160.000000 559.850000 1165.000000 560.150000 ;
        RECT 1160.000000 583.850000 1165.000000 584.150000 ;
        RECT 1160.000000 567.850000 1165.000000 568.150000 ;
        RECT 1160.000000 571.850000 1165.000000 572.150000 ;
        RECT 1160.000000 579.850000 1165.000000 580.150000 ;
        RECT 1160.000000 575.850000 1165.000000 576.150000 ;
        RECT 1160.000000 591.850000 1165.000000 592.150000 ;
        RECT 1160.000000 587.850000 1165.000000 588.150000 ;
        RECT 1160.000000 595.850000 1165.000000 596.150000 ;
        RECT 1160.000000 599.850000 1165.000000 600.150000 ;
        RECT 1160.000000 607.850000 1165.000000 608.150000 ;
        RECT 1160.000000 603.850000 1165.000000 604.150000 ;
        RECT 1160.000000 611.850000 1165.000000 612.150000 ;
        RECT 1160.000000 615.850000 1165.000000 616.150000 ;
        RECT 1160.000000 619.850000 1165.000000 620.150000 ;
        RECT 1160.000000 623.850000 1165.000000 624.150000 ;
        RECT 1160.000000 627.850000 1165.000000 628.150000 ;
        RECT 1160.000000 635.850000 1165.000000 636.150000 ;
        RECT 1160.000000 631.850000 1165.000000 632.150000 ;
        RECT 610.000000 659.850000 615.000000 660.150000 ;
        RECT 610.000000 663.850000 615.000000 664.150000 ;
        RECT 610.000000 667.850000 615.000000 668.150000 ;
        RECT 610.000000 671.850000 615.000000 672.150000 ;
        RECT 610.000000 675.850000 615.000000 676.150000 ;
        RECT 660.000000 663.850000 665.000000 664.150000 ;
        RECT 660.000000 659.850000 665.000000 660.150000 ;
        RECT 660.000000 667.850000 665.000000 668.150000 ;
        RECT 660.000000 671.850000 665.000000 672.150000 ;
        RECT 660.000000 675.850000 665.000000 676.150000 ;
        RECT 610.000000 683.850000 615.000000 684.150000 ;
        RECT 610.000000 679.850000 615.000000 680.150000 ;
        RECT 660.000000 683.850000 665.000000 684.150000 ;
        RECT 660.000000 679.850000 665.000000 680.150000 ;
        RECT 1160.000000 639.850000 1165.000000 640.150000 ;
        RECT 1160.000000 643.850000 1165.000000 644.150000 ;
        RECT 1160.000000 647.850000 1165.000000 648.150000 ;
        RECT 1160.000000 655.850000 1165.000000 656.150000 ;
        RECT 1160.000000 651.850000 1165.000000 652.150000 ;
        RECT 1160.000000 663.850000 1165.000000 664.150000 ;
        RECT 1160.000000 659.850000 1165.000000 660.150000 ;
        RECT 1160.000000 667.850000 1165.000000 668.150000 ;
        RECT 1160.000000 671.850000 1165.000000 672.150000 ;
        RECT 1160.000000 675.850000 1165.000000 676.150000 ;
        RECT 1160.000000 683.850000 1165.000000 684.150000 ;
        RECT 1160.000000 679.850000 1165.000000 680.150000 ;
      LAYER M3 ;
        RECT 60.000000 3.850000 65.000000 4.150000 ;
        RECT 60.000000 7.850000 65.000000 8.150000 ;
        RECT 110.000000 7.850000 115.000000 8.150000 ;
        RECT 110.000000 3.850000 115.000000 4.150000 ;
        RECT 160.000000 7.850000 165.000000 8.150000 ;
        RECT 160.000000 3.850000 165.000000 4.150000 ;
        RECT 210.000000 7.850000 215.000000 8.150000 ;
        RECT 210.000000 3.850000 215.000000 4.150000 ;
        RECT 260.000000 7.850000 265.000000 8.150000 ;
        RECT 260.000000 3.850000 265.000000 4.150000 ;
        RECT 310.000000 7.850000 315.000000 8.150000 ;
        RECT 310.000000 3.850000 315.000000 4.150000 ;
        RECT 360.000000 7.850000 365.000000 8.150000 ;
        RECT 360.000000 3.850000 365.000000 4.150000 ;
        RECT 410.000000 7.850000 415.000000 8.150000 ;
        RECT 410.000000 3.850000 415.000000 4.150000 ;
        RECT 460.000000 7.850000 465.000000 8.150000 ;
        RECT 460.000000 3.850000 465.000000 4.150000 ;
        RECT 510.000000 7.850000 515.000000 8.150000 ;
        RECT 510.000000 3.850000 515.000000 4.150000 ;
        RECT 560.000000 7.850000 565.000000 8.150000 ;
        RECT 560.000000 3.850000 565.000000 4.150000 ;
        RECT 18.000000 259.850000 28.000000 260.150000 ;
        RECT 18.000000 263.850000 28.000000 264.150000 ;
        RECT 18.000000 267.850000 28.000000 268.150000 ;
        RECT 60.000000 267.850000 65.000000 268.150000 ;
        RECT 60.000000 263.850000 65.000000 264.150000 ;
        RECT 60.000000 259.850000 65.000000 260.150000 ;
        RECT 110.000000 267.850000 115.000000 268.150000 ;
        RECT 110.000000 259.850000 115.000000 260.150000 ;
        RECT 110.000000 263.850000 115.000000 264.150000 ;
        RECT 18.000000 283.850000 28.000000 284.150000 ;
        RECT 18.000000 279.850000 28.000000 280.150000 ;
        RECT 18.000000 275.850000 28.000000 276.150000 ;
        RECT 18.000000 271.850000 28.000000 272.150000 ;
        RECT 18.000000 287.850000 28.000000 288.150000 ;
        RECT 18.000000 291.850000 28.000000 292.150000 ;
        RECT 18.000000 295.850000 28.000000 296.150000 ;
        RECT 18.000000 299.850000 28.000000 300.150000 ;
        RECT 18.000000 303.850000 28.000000 304.150000 ;
        RECT 60.000000 283.850000 65.000000 284.150000 ;
        RECT 60.000000 279.850000 65.000000 280.150000 ;
        RECT 60.000000 275.850000 65.000000 276.150000 ;
        RECT 60.000000 271.850000 65.000000 272.150000 ;
        RECT 60.000000 287.850000 65.000000 288.150000 ;
        RECT 60.000000 291.850000 65.000000 292.150000 ;
        RECT 60.000000 295.850000 65.000000 296.150000 ;
        RECT 60.000000 299.850000 65.000000 300.150000 ;
        RECT 60.000000 303.850000 65.000000 304.150000 ;
        RECT 18.000000 307.850000 28.000000 308.150000 ;
        RECT 18.000000 311.850000 28.000000 312.150000 ;
        RECT 18.000000 315.850000 28.000000 316.150000 ;
        RECT 18.000000 319.850000 28.000000 320.150000 ;
        RECT 18.000000 323.850000 28.000000 324.150000 ;
        RECT 18.000000 339.850000 28.000000 340.150000 ;
        RECT 18.000000 335.850000 28.000000 336.150000 ;
        RECT 18.000000 331.850000 28.000000 332.150000 ;
        RECT 18.000000 327.850000 28.000000 328.150000 ;
        RECT 60.000000 307.850000 65.000000 308.150000 ;
        RECT 60.000000 311.850000 65.000000 312.150000 ;
        RECT 60.000000 315.850000 65.000000 316.150000 ;
        RECT 60.000000 319.850000 65.000000 320.150000 ;
        RECT 60.000000 323.850000 65.000000 324.150000 ;
        RECT 60.000000 339.850000 65.000000 340.150000 ;
        RECT 60.000000 335.850000 65.000000 336.150000 ;
        RECT 60.000000 331.850000 65.000000 332.150000 ;
        RECT 60.000000 327.850000 65.000000 328.150000 ;
        RECT 110.000000 271.850000 115.000000 272.150000 ;
        RECT 110.000000 275.850000 115.000000 276.150000 ;
        RECT 110.000000 279.850000 115.000000 280.150000 ;
        RECT 110.000000 283.850000 115.000000 284.150000 ;
        RECT 110.000000 287.850000 115.000000 288.150000 ;
        RECT 110.000000 291.850000 115.000000 292.150000 ;
        RECT 110.000000 295.850000 115.000000 296.150000 ;
        RECT 110.000000 299.850000 115.000000 300.150000 ;
        RECT 110.000000 303.850000 115.000000 304.150000 ;
        RECT 110.000000 311.850000 115.000000 312.150000 ;
        RECT 110.000000 307.850000 115.000000 308.150000 ;
        RECT 110.000000 323.850000 115.000000 324.150000 ;
        RECT 110.000000 319.850000 115.000000 320.150000 ;
        RECT 110.000000 315.850000 115.000000 316.150000 ;
        RECT 110.000000 339.850000 115.000000 340.150000 ;
        RECT 110.000000 335.850000 115.000000 336.150000 ;
        RECT 110.000000 331.850000 115.000000 332.150000 ;
        RECT 110.000000 327.850000 115.000000 328.150000 ;
        RECT 160.000000 259.850000 165.000000 260.150000 ;
        RECT 160.000000 263.850000 165.000000 264.150000 ;
        RECT 160.000000 267.850000 165.000000 268.150000 ;
        RECT 210.000000 267.850000 215.000000 268.150000 ;
        RECT 210.000000 263.850000 215.000000 264.150000 ;
        RECT 210.000000 259.850000 215.000000 260.150000 ;
        RECT 260.000000 267.850000 265.000000 268.150000 ;
        RECT 260.000000 259.850000 265.000000 260.150000 ;
        RECT 260.000000 263.850000 265.000000 264.150000 ;
        RECT 160.000000 275.850000 165.000000 276.150000 ;
        RECT 160.000000 271.850000 165.000000 272.150000 ;
        RECT 160.000000 283.850000 165.000000 284.150000 ;
        RECT 160.000000 279.850000 165.000000 280.150000 ;
        RECT 160.000000 287.850000 165.000000 288.150000 ;
        RECT 160.000000 291.850000 165.000000 292.150000 ;
        RECT 160.000000 295.850000 165.000000 296.150000 ;
        RECT 160.000000 299.850000 165.000000 300.150000 ;
        RECT 160.000000 303.850000 165.000000 304.150000 ;
        RECT 210.000000 283.850000 215.000000 284.150000 ;
        RECT 210.000000 279.850000 215.000000 280.150000 ;
        RECT 210.000000 275.850000 215.000000 276.150000 ;
        RECT 210.000000 271.850000 215.000000 272.150000 ;
        RECT 210.000000 287.850000 215.000000 288.150000 ;
        RECT 210.000000 291.850000 215.000000 292.150000 ;
        RECT 210.000000 295.850000 215.000000 296.150000 ;
        RECT 210.000000 299.850000 215.000000 300.150000 ;
        RECT 210.000000 303.850000 215.000000 304.150000 ;
        RECT 160.000000 311.850000 165.000000 312.150000 ;
        RECT 160.000000 307.850000 165.000000 308.150000 ;
        RECT 160.000000 315.850000 165.000000 316.150000 ;
        RECT 160.000000 319.850000 165.000000 320.150000 ;
        RECT 160.000000 323.850000 165.000000 324.150000 ;
        RECT 160.000000 331.850000 165.000000 332.150000 ;
        RECT 160.000000 327.850000 165.000000 328.150000 ;
        RECT 160.000000 335.850000 165.000000 336.150000 ;
        RECT 160.000000 339.850000 165.000000 340.150000 ;
        RECT 210.000000 307.850000 215.000000 308.150000 ;
        RECT 210.000000 311.850000 215.000000 312.150000 ;
        RECT 210.000000 315.850000 215.000000 316.150000 ;
        RECT 210.000000 323.850000 215.000000 324.150000 ;
        RECT 210.000000 319.850000 215.000000 320.150000 ;
        RECT 210.000000 327.850000 215.000000 328.150000 ;
        RECT 210.000000 331.850000 215.000000 332.150000 ;
        RECT 210.000000 335.850000 215.000000 336.150000 ;
        RECT 210.000000 339.850000 215.000000 340.150000 ;
        RECT 260.000000 271.850000 265.000000 272.150000 ;
        RECT 260.000000 275.850000 265.000000 276.150000 ;
        RECT 260.000000 279.850000 265.000000 280.150000 ;
        RECT 260.000000 283.850000 265.000000 284.150000 ;
        RECT 260.000000 291.850000 265.000000 292.150000 ;
        RECT 260.000000 287.850000 265.000000 288.150000 ;
        RECT 260.000000 295.850000 265.000000 296.150000 ;
        RECT 260.000000 303.850000 265.000000 304.150000 ;
        RECT 260.000000 299.850000 265.000000 300.150000 ;
        RECT 260.000000 307.850000 265.000000 308.150000 ;
        RECT 260.000000 311.850000 265.000000 312.150000 ;
        RECT 260.000000 315.850000 265.000000 316.150000 ;
        RECT 260.000000 319.850000 265.000000 320.150000 ;
        RECT 260.000000 323.850000 265.000000 324.150000 ;
        RECT 260.000000 327.850000 265.000000 328.150000 ;
        RECT 260.000000 331.850000 265.000000 332.150000 ;
        RECT 260.000000 335.850000 265.000000 336.150000 ;
        RECT 260.000000 339.850000 265.000000 340.150000 ;
        RECT 310.000000 259.850000 315.000000 260.150000 ;
        RECT 310.000000 263.850000 315.000000 264.150000 ;
        RECT 310.000000 267.850000 315.000000 268.150000 ;
        RECT 360.000000 267.850000 365.000000 268.150000 ;
        RECT 360.000000 263.850000 365.000000 264.150000 ;
        RECT 360.000000 259.850000 365.000000 260.150000 ;
        RECT 410.000000 259.850000 415.000000 260.150000 ;
        RECT 410.000000 263.850000 415.000000 264.150000 ;
        RECT 410.000000 267.850000 415.000000 268.150000 ;
        RECT 310.000000 275.850000 315.000000 276.150000 ;
        RECT 310.000000 271.850000 315.000000 272.150000 ;
        RECT 310.000000 283.850000 315.000000 284.150000 ;
        RECT 310.000000 279.850000 315.000000 280.150000 ;
        RECT 310.000000 291.850000 315.000000 292.150000 ;
        RECT 310.000000 287.850000 315.000000 288.150000 ;
        RECT 310.000000 295.850000 315.000000 296.150000 ;
        RECT 310.000000 303.850000 315.000000 304.150000 ;
        RECT 310.000000 299.850000 315.000000 300.150000 ;
        RECT 360.000000 283.850000 365.000000 284.150000 ;
        RECT 360.000000 279.850000 365.000000 280.150000 ;
        RECT 360.000000 275.850000 365.000000 276.150000 ;
        RECT 360.000000 271.850000 365.000000 272.150000 ;
        RECT 360.000000 287.850000 365.000000 288.150000 ;
        RECT 360.000000 291.850000 365.000000 292.150000 ;
        RECT 360.000000 295.850000 365.000000 296.150000 ;
        RECT 360.000000 299.850000 365.000000 300.150000 ;
        RECT 360.000000 303.850000 365.000000 304.150000 ;
        RECT 310.000000 311.850000 315.000000 312.150000 ;
        RECT 310.000000 307.850000 315.000000 308.150000 ;
        RECT 310.000000 315.850000 315.000000 316.150000 ;
        RECT 310.000000 323.850000 315.000000 324.150000 ;
        RECT 310.000000 319.850000 315.000000 320.150000 ;
        RECT 310.000000 327.850000 315.000000 328.150000 ;
        RECT 310.000000 331.850000 315.000000 332.150000 ;
        RECT 310.000000 335.850000 315.000000 336.150000 ;
        RECT 310.000000 339.850000 315.000000 340.150000 ;
        RECT 360.000000 307.850000 365.000000 308.150000 ;
        RECT 360.000000 311.850000 365.000000 312.150000 ;
        RECT 360.000000 315.850000 365.000000 316.150000 ;
        RECT 360.000000 319.850000 365.000000 320.150000 ;
        RECT 360.000000 323.850000 365.000000 324.150000 ;
        RECT 360.000000 339.850000 365.000000 340.150000 ;
        RECT 360.000000 335.850000 365.000000 336.150000 ;
        RECT 360.000000 331.850000 365.000000 332.150000 ;
        RECT 360.000000 327.850000 365.000000 328.150000 ;
        RECT 410.000000 271.850000 415.000000 272.150000 ;
        RECT 410.000000 275.850000 415.000000 276.150000 ;
        RECT 410.000000 279.850000 415.000000 280.150000 ;
        RECT 410.000000 283.850000 415.000000 284.150000 ;
        RECT 410.000000 291.850000 415.000000 292.150000 ;
        RECT 410.000000 287.850000 415.000000 288.150000 ;
        RECT 410.000000 295.850000 415.000000 296.150000 ;
        RECT 410.000000 299.850000 415.000000 300.150000 ;
        RECT 410.000000 303.850000 415.000000 304.150000 ;
        RECT 410.000000 307.850000 415.000000 308.150000 ;
        RECT 410.000000 311.850000 415.000000 312.150000 ;
        RECT 410.000000 315.850000 415.000000 316.150000 ;
        RECT 410.000000 319.850000 415.000000 320.150000 ;
        RECT 410.000000 323.850000 415.000000 324.150000 ;
        RECT 410.000000 327.850000 415.000000 328.150000 ;
        RECT 410.000000 331.850000 415.000000 332.150000 ;
        RECT 410.000000 339.850000 415.000000 340.150000 ;
        RECT 410.000000 335.850000 415.000000 336.150000 ;
        RECT 460.000000 259.850000 465.000000 260.150000 ;
        RECT 460.000000 263.850000 465.000000 264.150000 ;
        RECT 460.000000 267.850000 465.000000 268.150000 ;
        RECT 510.000000 259.850000 515.000000 260.150000 ;
        RECT 510.000000 263.850000 515.000000 264.150000 ;
        RECT 510.000000 267.850000 515.000000 268.150000 ;
        RECT 560.000000 263.850000 565.000000 264.150000 ;
        RECT 560.000000 259.850000 565.000000 260.150000 ;
        RECT 560.000000 267.850000 565.000000 268.150000 ;
        RECT 460.000000 283.850000 465.000000 284.150000 ;
        RECT 460.000000 279.850000 465.000000 280.150000 ;
        RECT 460.000000 275.850000 465.000000 276.150000 ;
        RECT 460.000000 271.850000 465.000000 272.150000 ;
        RECT 460.000000 295.850000 465.000000 296.150000 ;
        RECT 460.000000 291.850000 465.000000 292.150000 ;
        RECT 460.000000 287.850000 465.000000 288.150000 ;
        RECT 460.000000 301.230000 465.000000 302.230000 ;
        RECT 510.000000 271.850000 515.000000 272.150000 ;
        RECT 510.000000 275.850000 515.000000 276.150000 ;
        RECT 510.000000 279.850000 515.000000 280.150000 ;
        RECT 510.000000 283.850000 515.000000 284.150000 ;
        RECT 510.000000 291.850000 515.000000 292.150000 ;
        RECT 510.000000 287.850000 515.000000 288.150000 ;
        RECT 510.000000 295.850000 515.000000 296.150000 ;
        RECT 510.000000 299.850000 515.000000 300.150000 ;
        RECT 510.000000 303.850000 515.000000 304.150000 ;
        RECT 460.000000 319.850000 465.000000 320.150000 ;
        RECT 460.000000 323.850000 465.000000 324.150000 ;
        RECT 460.000000 339.850000 465.000000 340.150000 ;
        RECT 460.000000 335.850000 465.000000 336.150000 ;
        RECT 460.000000 331.850000 465.000000 332.150000 ;
        RECT 460.000000 327.850000 465.000000 328.150000 ;
        RECT 510.000000 311.850000 515.000000 312.150000 ;
        RECT 510.000000 307.850000 515.000000 308.150000 ;
        RECT 510.000000 315.850000 515.000000 316.150000 ;
        RECT 510.000000 323.850000 515.000000 324.150000 ;
        RECT 510.000000 319.850000 515.000000 320.150000 ;
        RECT 510.000000 331.850000 515.000000 332.150000 ;
        RECT 510.000000 327.850000 515.000000 328.150000 ;
        RECT 510.000000 335.850000 515.000000 336.150000 ;
        RECT 510.000000 339.850000 515.000000 340.150000 ;
        RECT 560.000000 283.850000 565.000000 284.150000 ;
        RECT 560.000000 279.850000 565.000000 280.150000 ;
        RECT 560.000000 275.850000 565.000000 276.150000 ;
        RECT 560.000000 271.850000 565.000000 272.150000 ;
        RECT 560.000000 287.850000 565.000000 288.150000 ;
        RECT 560.000000 291.850000 565.000000 292.150000 ;
        RECT 560.000000 295.850000 565.000000 296.150000 ;
        RECT 560.000000 299.850000 565.000000 300.150000 ;
        RECT 560.000000 303.850000 565.000000 304.150000 ;
        RECT 560.000000 323.850000 565.000000 324.150000 ;
        RECT 560.000000 319.850000 565.000000 320.150000 ;
        RECT 560.000000 315.850000 565.000000 316.150000 ;
        RECT 560.000000 311.850000 565.000000 312.150000 ;
        RECT 560.000000 307.850000 565.000000 308.150000 ;
        RECT 560.000000 339.850000 565.000000 340.150000 ;
        RECT 560.000000 335.850000 565.000000 336.150000 ;
        RECT 560.000000 331.850000 565.000000 332.150000 ;
        RECT 560.000000 327.850000 565.000000 328.150000 ;
        RECT 610.000000 7.850000 615.000000 8.150000 ;
        RECT 610.000000 3.850000 615.000000 4.150000 ;
        RECT 660.000000 7.850000 665.000000 8.150000 ;
        RECT 660.000000 3.850000 665.000000 4.150000 ;
        RECT 710.000000 7.850000 715.000000 8.150000 ;
        RECT 710.000000 3.850000 715.000000 4.150000 ;
        RECT 760.000000 7.850000 765.000000 8.150000 ;
        RECT 760.000000 3.850000 765.000000 4.150000 ;
        RECT 810.000000 7.850000 815.000000 8.150000 ;
        RECT 810.000000 3.850000 815.000000 4.150000 ;
        RECT 860.000000 7.850000 865.000000 8.150000 ;
        RECT 860.000000 3.850000 865.000000 4.150000 ;
        RECT 960.000000 7.850000 965.000000 8.150000 ;
        RECT 960.000000 3.850000 965.000000 4.150000 ;
        RECT 910.000000 7.850000 915.000000 8.150000 ;
        RECT 910.000000 3.850000 915.000000 4.150000 ;
        RECT 1010.000000 7.850000 1015.000000 8.150000 ;
        RECT 1010.000000 3.850000 1015.000000 4.150000 ;
        RECT 1110.000000 7.850000 1115.000000 8.150000 ;
        RECT 1110.000000 3.850000 1115.000000 4.150000 ;
        RECT 1060.000000 7.850000 1065.000000 8.150000 ;
        RECT 1060.000000 3.850000 1065.000000 4.150000 ;
        RECT 1160.000000 3.850000 1165.000000 4.150000 ;
        RECT 1160.000000 7.850000 1165.000000 8.150000 ;
        RECT 1158.000000 27.850000 1168.000000 28.150000 ;
        RECT 1158.000000 23.850000 1168.000000 24.150000 ;
        RECT 1158.000000 19.850000 1168.000000 20.150000 ;
        RECT 1160.000000 15.850000 1165.000000 16.150000 ;
        RECT 1160.000000 11.850000 1165.000000 12.150000 ;
        RECT 1158.000000 31.850000 1168.000000 32.150000 ;
        RECT 1158.000000 35.850000 1168.000000 36.150000 ;
        RECT 1158.000000 43.850000 1168.000000 44.150000 ;
        RECT 1158.000000 39.850000 1168.000000 40.150000 ;
        RECT 610.000000 267.850000 615.000000 268.150000 ;
        RECT 610.000000 263.850000 615.000000 264.150000 ;
        RECT 610.000000 259.850000 615.000000 260.150000 ;
        RECT 660.000000 259.850000 665.000000 260.150000 ;
        RECT 660.000000 263.850000 665.000000 264.150000 ;
        RECT 660.000000 267.850000 665.000000 268.150000 ;
        RECT 710.000000 267.850000 715.000000 268.150000 ;
        RECT 710.000000 259.850000 715.000000 260.150000 ;
        RECT 710.000000 263.850000 715.000000 264.150000 ;
        RECT 610.000000 283.850000 615.000000 284.150000 ;
        RECT 610.000000 279.850000 615.000000 280.150000 ;
        RECT 610.000000 275.850000 615.000000 276.150000 ;
        RECT 610.000000 271.850000 615.000000 272.150000 ;
        RECT 610.000000 287.850000 615.000000 288.150000 ;
        RECT 610.000000 291.850000 615.000000 292.150000 ;
        RECT 610.000000 295.850000 615.000000 296.150000 ;
        RECT 610.000000 299.850000 615.000000 300.150000 ;
        RECT 610.000000 303.850000 615.000000 304.150000 ;
        RECT 660.000000 275.850000 665.000000 276.150000 ;
        RECT 660.000000 271.850000 665.000000 272.150000 ;
        RECT 660.000000 283.850000 665.000000 284.150000 ;
        RECT 660.000000 279.850000 665.000000 280.150000 ;
        RECT 660.000000 287.850000 665.000000 288.150000 ;
        RECT 660.000000 291.850000 665.000000 292.150000 ;
        RECT 660.000000 295.850000 665.000000 296.150000 ;
        RECT 660.000000 303.850000 665.000000 304.150000 ;
        RECT 660.000000 299.850000 665.000000 300.150000 ;
        RECT 610.000000 307.850000 615.000000 308.150000 ;
        RECT 610.000000 311.850000 615.000000 312.150000 ;
        RECT 610.000000 315.850000 615.000000 316.150000 ;
        RECT 610.000000 319.850000 615.000000 320.150000 ;
        RECT 610.000000 323.850000 615.000000 324.150000 ;
        RECT 610.000000 339.850000 615.000000 340.150000 ;
        RECT 610.000000 335.850000 615.000000 336.150000 ;
        RECT 610.000000 331.850000 615.000000 332.150000 ;
        RECT 610.000000 327.850000 615.000000 328.150000 ;
        RECT 660.000000 311.850000 665.000000 312.150000 ;
        RECT 660.000000 307.850000 665.000000 308.150000 ;
        RECT 660.000000 315.850000 665.000000 316.150000 ;
        RECT 660.000000 319.850000 665.000000 320.150000 ;
        RECT 660.000000 323.850000 665.000000 324.150000 ;
        RECT 660.000000 331.850000 665.000000 332.150000 ;
        RECT 660.000000 327.850000 665.000000 328.150000 ;
        RECT 660.000000 335.850000 665.000000 336.150000 ;
        RECT 660.000000 339.850000 665.000000 340.150000 ;
        RECT 710.000000 271.850000 715.000000 272.150000 ;
        RECT 710.000000 275.850000 715.000000 276.150000 ;
        RECT 710.000000 279.850000 715.000000 280.150000 ;
        RECT 710.000000 283.850000 715.000000 284.150000 ;
        RECT 710.000000 287.850000 715.000000 288.150000 ;
        RECT 710.000000 291.850000 715.000000 292.150000 ;
        RECT 710.000000 295.850000 715.000000 296.150000 ;
        RECT 710.000000 299.850000 715.000000 300.150000 ;
        RECT 710.000000 303.850000 715.000000 304.150000 ;
        RECT 710.000000 323.850000 715.000000 324.150000 ;
        RECT 710.000000 319.850000 715.000000 320.150000 ;
        RECT 710.000000 315.850000 715.000000 316.150000 ;
        RECT 710.000000 311.850000 715.000000 312.150000 ;
        RECT 710.000000 307.850000 715.000000 308.150000 ;
        RECT 710.000000 339.850000 715.000000 340.150000 ;
        RECT 710.000000 335.850000 715.000000 336.150000 ;
        RECT 710.000000 331.850000 715.000000 332.150000 ;
        RECT 710.000000 327.850000 715.000000 328.150000 ;
        RECT 760.000000 267.850000 765.000000 268.150000 ;
        RECT 760.000000 263.850000 765.000000 264.150000 ;
        RECT 760.000000 259.850000 765.000000 260.150000 ;
        RECT 810.000000 259.850000 815.000000 260.150000 ;
        RECT 810.000000 263.850000 815.000000 264.150000 ;
        RECT 810.000000 267.850000 815.000000 268.150000 ;
        RECT 860.000000 267.850000 865.000000 268.150000 ;
        RECT 860.000000 259.850000 865.000000 260.150000 ;
        RECT 860.000000 263.850000 865.000000 264.150000 ;
        RECT 760.000000 283.850000 765.000000 284.150000 ;
        RECT 760.000000 279.850000 765.000000 280.150000 ;
        RECT 760.000000 275.850000 765.000000 276.150000 ;
        RECT 760.000000 271.850000 765.000000 272.150000 ;
        RECT 760.000000 287.850000 765.000000 288.150000 ;
        RECT 760.000000 291.850000 765.000000 292.150000 ;
        RECT 760.000000 295.850000 765.000000 296.150000 ;
        RECT 760.000000 299.850000 765.000000 300.150000 ;
        RECT 760.000000 303.850000 765.000000 304.150000 ;
        RECT 810.000000 275.850000 815.000000 276.150000 ;
        RECT 810.000000 271.850000 815.000000 272.150000 ;
        RECT 810.000000 283.850000 815.000000 284.150000 ;
        RECT 810.000000 279.850000 815.000000 280.150000 ;
        RECT 810.000000 287.850000 815.000000 288.150000 ;
        RECT 810.000000 291.850000 815.000000 292.150000 ;
        RECT 810.000000 295.850000 815.000000 296.150000 ;
        RECT 810.000000 303.850000 815.000000 304.150000 ;
        RECT 810.000000 299.850000 815.000000 300.150000 ;
        RECT 760.000000 307.850000 765.000000 308.150000 ;
        RECT 760.000000 311.850000 765.000000 312.150000 ;
        RECT 760.000000 315.850000 765.000000 316.150000 ;
        RECT 760.000000 319.850000 765.000000 320.150000 ;
        RECT 760.000000 323.850000 765.000000 324.150000 ;
        RECT 760.000000 339.850000 765.000000 340.150000 ;
        RECT 760.000000 335.850000 765.000000 336.150000 ;
        RECT 760.000000 331.850000 765.000000 332.150000 ;
        RECT 760.000000 327.850000 765.000000 328.150000 ;
        RECT 810.000000 311.850000 815.000000 312.150000 ;
        RECT 810.000000 307.850000 815.000000 308.150000 ;
        RECT 810.000000 315.850000 815.000000 316.150000 ;
        RECT 810.000000 319.850000 815.000000 320.150000 ;
        RECT 810.000000 323.850000 815.000000 324.150000 ;
        RECT 810.000000 331.850000 815.000000 332.150000 ;
        RECT 810.000000 327.850000 815.000000 328.150000 ;
        RECT 810.000000 335.850000 815.000000 336.150000 ;
        RECT 810.000000 339.850000 815.000000 340.150000 ;
        RECT 860.000000 271.850000 865.000000 272.150000 ;
        RECT 860.000000 275.850000 865.000000 276.150000 ;
        RECT 860.000000 279.850000 865.000000 280.150000 ;
        RECT 860.000000 283.850000 865.000000 284.150000 ;
        RECT 860.000000 287.850000 865.000000 288.150000 ;
        RECT 860.000000 291.850000 865.000000 292.150000 ;
        RECT 860.000000 295.850000 865.000000 296.150000 ;
        RECT 860.000000 299.850000 865.000000 300.150000 ;
        RECT 860.000000 303.850000 865.000000 304.150000 ;
        RECT 860.000000 323.850000 865.000000 324.150000 ;
        RECT 860.000000 319.850000 865.000000 320.150000 ;
        RECT 860.000000 315.850000 865.000000 316.150000 ;
        RECT 860.000000 311.850000 865.000000 312.150000 ;
        RECT 860.000000 307.850000 865.000000 308.150000 ;
        RECT 860.000000 339.850000 865.000000 340.150000 ;
        RECT 860.000000 335.850000 865.000000 336.150000 ;
        RECT 860.000000 331.850000 865.000000 332.150000 ;
        RECT 860.000000 327.850000 865.000000 328.150000 ;
        RECT 1158.000000 47.850000 1168.000000 48.150000 ;
        RECT 1158.000000 51.850000 1168.000000 52.150000 ;
        RECT 1158.000000 63.850000 1168.000000 64.150000 ;
        RECT 1158.000000 55.850000 1168.000000 56.150000 ;
        RECT 1158.000000 59.850000 1168.000000 60.150000 ;
        RECT 1158.000000 67.850000 1168.000000 68.150000 ;
        RECT 1158.000000 71.850000 1168.000000 72.150000 ;
        RECT 1158.000000 79.850000 1168.000000 80.150000 ;
        RECT 1158.000000 75.850000 1168.000000 76.150000 ;
        RECT 1158.000000 83.850000 1168.000000 84.150000 ;
        RECT 1158.000000 87.850000 1168.000000 88.150000 ;
        RECT 1158.000000 91.850000 1168.000000 92.150000 ;
        RECT 1158.000000 99.850000 1168.000000 100.150000 ;
        RECT 1158.000000 95.850000 1168.000000 96.150000 ;
        RECT 1158.000000 103.850000 1168.000000 104.150000 ;
        RECT 1158.000000 107.850000 1168.000000 108.150000 ;
        RECT 1158.000000 119.850000 1168.000000 120.150000 ;
        RECT 1158.000000 115.850000 1168.000000 116.150000 ;
        RECT 1158.000000 111.850000 1168.000000 112.150000 ;
        RECT 1158.000000 123.850000 1168.000000 124.150000 ;
        RECT 1158.000000 127.850000 1168.000000 128.150000 ;
        RECT 1158.000000 135.850000 1168.000000 136.150000 ;
        RECT 1158.000000 131.850000 1168.000000 132.150000 ;
        RECT 1158.000000 139.850000 1168.000000 140.150000 ;
        RECT 1158.000000 143.850000 1168.000000 144.150000 ;
        RECT 1158.000000 147.850000 1168.000000 148.150000 ;
        RECT 1158.000000 155.850000 1168.000000 156.150000 ;
        RECT 1158.000000 151.850000 1168.000000 152.150000 ;
        RECT 1158.000000 159.850000 1168.000000 160.150000 ;
        RECT 1158.000000 163.850000 1168.000000 164.150000 ;
        RECT 1158.000000 175.850000 1168.000000 176.150000 ;
        RECT 1158.000000 171.850000 1168.000000 172.150000 ;
        RECT 1158.000000 167.850000 1168.000000 168.150000 ;
        RECT 1158.000000 179.850000 1168.000000 180.150000 ;
        RECT 1158.000000 183.850000 1168.000000 184.150000 ;
        RECT 1158.000000 191.850000 1168.000000 192.150000 ;
        RECT 1158.000000 187.850000 1168.000000 188.150000 ;
        RECT 960.000000 267.850000 965.000000 268.150000 ;
        RECT 960.000000 263.850000 965.000000 264.150000 ;
        RECT 960.000000 259.850000 965.000000 260.150000 ;
        RECT 910.000000 267.850000 915.000000 268.150000 ;
        RECT 910.000000 263.850000 915.000000 264.150000 ;
        RECT 910.000000 259.850000 915.000000 260.150000 ;
        RECT 1010.000000 259.850000 1015.000000 260.150000 ;
        RECT 1010.000000 263.850000 1015.000000 264.150000 ;
        RECT 1010.000000 267.850000 1015.000000 268.150000 ;
        RECT 960.000000 283.850000 965.000000 284.150000 ;
        RECT 960.000000 279.850000 965.000000 280.150000 ;
        RECT 960.000000 275.850000 965.000000 276.150000 ;
        RECT 960.000000 271.850000 965.000000 272.150000 ;
        RECT 960.000000 287.850000 965.000000 288.150000 ;
        RECT 960.000000 291.850000 965.000000 292.150000 ;
        RECT 960.000000 295.850000 965.000000 296.150000 ;
        RECT 960.000000 299.850000 965.000000 300.150000 ;
        RECT 960.000000 303.850000 965.000000 304.150000 ;
        RECT 960.000000 311.850000 965.000000 312.150000 ;
        RECT 960.000000 307.850000 965.000000 308.150000 ;
        RECT 960.000000 323.850000 965.000000 324.150000 ;
        RECT 960.000000 319.850000 965.000000 320.150000 ;
        RECT 960.000000 315.850000 965.000000 316.150000 ;
        RECT 960.000000 339.850000 965.000000 340.150000 ;
        RECT 960.000000 335.850000 965.000000 336.150000 ;
        RECT 960.000000 331.850000 965.000000 332.150000 ;
        RECT 960.000000 327.850000 965.000000 328.150000 ;
        RECT 910.000000 283.850000 915.000000 284.150000 ;
        RECT 910.000000 279.850000 915.000000 280.150000 ;
        RECT 910.000000 275.850000 915.000000 276.150000 ;
        RECT 910.000000 271.850000 915.000000 272.150000 ;
        RECT 910.000000 287.850000 915.000000 288.150000 ;
        RECT 910.000000 291.850000 915.000000 292.150000 ;
        RECT 910.000000 295.850000 915.000000 296.150000 ;
        RECT 910.000000 299.850000 915.000000 300.150000 ;
        RECT 910.000000 303.850000 915.000000 304.150000 ;
        RECT 910.000000 307.850000 915.000000 308.150000 ;
        RECT 910.000000 311.850000 915.000000 312.150000 ;
        RECT 910.000000 315.850000 915.000000 316.150000 ;
        RECT 910.000000 319.850000 915.000000 320.150000 ;
        RECT 910.000000 323.850000 915.000000 324.150000 ;
        RECT 910.000000 339.850000 915.000000 340.150000 ;
        RECT 910.000000 335.850000 915.000000 336.150000 ;
        RECT 910.000000 331.850000 915.000000 332.150000 ;
        RECT 910.000000 327.850000 915.000000 328.150000 ;
        RECT 1010.000000 275.850000 1015.000000 276.150000 ;
        RECT 1010.000000 271.850000 1015.000000 272.150000 ;
        RECT 1010.000000 283.850000 1015.000000 284.150000 ;
        RECT 1010.000000 279.850000 1015.000000 280.150000 ;
        RECT 1010.000000 287.850000 1015.000000 288.150000 ;
        RECT 1010.000000 291.850000 1015.000000 292.150000 ;
        RECT 1010.000000 295.850000 1015.000000 296.150000 ;
        RECT 1010.000000 303.850000 1015.000000 304.150000 ;
        RECT 1010.000000 299.850000 1015.000000 300.150000 ;
        RECT 1010.000000 311.850000 1015.000000 312.150000 ;
        RECT 1010.000000 307.850000 1015.000000 308.150000 ;
        RECT 1010.000000 315.850000 1015.000000 316.150000 ;
        RECT 1010.000000 319.850000 1015.000000 320.150000 ;
        RECT 1010.000000 323.850000 1015.000000 324.150000 ;
        RECT 1010.000000 331.850000 1015.000000 332.150000 ;
        RECT 1010.000000 327.850000 1015.000000 328.150000 ;
        RECT 1010.000000 335.850000 1015.000000 336.150000 ;
        RECT 1010.000000 339.850000 1015.000000 340.150000 ;
        RECT 1110.000000 267.850000 1115.000000 268.150000 ;
        RECT 1110.000000 263.850000 1115.000000 264.150000 ;
        RECT 1110.000000 259.850000 1115.000000 260.150000 ;
        RECT 1060.000000 267.850000 1065.000000 268.150000 ;
        RECT 1060.000000 263.850000 1065.000000 264.150000 ;
        RECT 1060.000000 259.850000 1065.000000 260.150000 ;
        RECT 1158.000000 203.850000 1168.000000 204.150000 ;
        RECT 1158.000000 195.850000 1168.000000 196.150000 ;
        RECT 1158.000000 199.850000 1168.000000 200.150000 ;
        RECT 1158.000000 211.850000 1168.000000 212.150000 ;
        RECT 1158.000000 207.850000 1168.000000 208.150000 ;
        RECT 1158.000000 215.850000 1168.000000 216.150000 ;
        RECT 1158.000000 219.850000 1168.000000 220.150000 ;
        RECT 1158.000000 227.850000 1168.000000 228.150000 ;
        RECT 1158.000000 223.850000 1168.000000 224.150000 ;
        RECT 1158.000000 231.850000 1168.000000 232.150000 ;
        RECT 1158.000000 235.850000 1168.000000 236.150000 ;
        RECT 1158.000000 239.850000 1168.000000 240.150000 ;
        RECT 1158.000000 247.850000 1168.000000 248.150000 ;
        RECT 1158.000000 243.850000 1168.000000 244.150000 ;
        RECT 1158.000000 251.850000 1168.000000 252.150000 ;
        RECT 1158.000000 255.850000 1168.000000 256.150000 ;
        RECT 1158.000000 267.850000 1168.000000 268.150000 ;
        RECT 1158.000000 259.850000 1168.000000 260.150000 ;
        RECT 1158.000000 263.850000 1168.000000 264.150000 ;
        RECT 1110.000000 283.850000 1115.000000 284.150000 ;
        RECT 1110.000000 279.850000 1115.000000 280.150000 ;
        RECT 1110.000000 275.850000 1115.000000 276.150000 ;
        RECT 1110.000000 271.850000 1115.000000 272.150000 ;
        RECT 1110.000000 287.850000 1115.000000 288.150000 ;
        RECT 1110.000000 291.850000 1115.000000 292.150000 ;
        RECT 1110.000000 295.850000 1115.000000 296.150000 ;
        RECT 1110.000000 299.850000 1115.000000 300.150000 ;
        RECT 1110.000000 303.850000 1115.000000 304.150000 ;
        RECT 1110.000000 311.850000 1115.000000 312.150000 ;
        RECT 1110.000000 307.850000 1115.000000 308.150000 ;
        RECT 1110.000000 323.850000 1115.000000 324.150000 ;
        RECT 1110.000000 319.850000 1115.000000 320.150000 ;
        RECT 1110.000000 315.850000 1115.000000 316.150000 ;
        RECT 1110.000000 339.850000 1115.000000 340.150000 ;
        RECT 1110.000000 335.850000 1115.000000 336.150000 ;
        RECT 1110.000000 331.850000 1115.000000 332.150000 ;
        RECT 1110.000000 327.850000 1115.000000 328.150000 ;
        RECT 1060.000000 283.850000 1065.000000 284.150000 ;
        RECT 1060.000000 279.850000 1065.000000 280.150000 ;
        RECT 1060.000000 275.850000 1065.000000 276.150000 ;
        RECT 1060.000000 271.850000 1065.000000 272.150000 ;
        RECT 1060.000000 287.850000 1065.000000 288.150000 ;
        RECT 1060.000000 291.850000 1065.000000 292.150000 ;
        RECT 1060.000000 295.850000 1065.000000 296.150000 ;
        RECT 1060.000000 299.850000 1065.000000 300.150000 ;
        RECT 1060.000000 303.850000 1065.000000 304.150000 ;
        RECT 1060.000000 307.850000 1065.000000 308.150000 ;
        RECT 1060.000000 311.850000 1065.000000 312.150000 ;
        RECT 1060.000000 315.850000 1065.000000 316.150000 ;
        RECT 1060.000000 319.850000 1065.000000 320.150000 ;
        RECT 1060.000000 323.850000 1065.000000 324.150000 ;
        RECT 1060.000000 339.850000 1065.000000 340.150000 ;
        RECT 1060.000000 335.850000 1065.000000 336.150000 ;
        RECT 1060.000000 331.850000 1065.000000 332.150000 ;
        RECT 1060.000000 327.850000 1065.000000 328.150000 ;
        RECT 1158.000000 283.850000 1168.000000 284.150000 ;
        RECT 1158.000000 279.850000 1168.000000 280.150000 ;
        RECT 1158.000000 275.850000 1168.000000 276.150000 ;
        RECT 1158.000000 271.850000 1168.000000 272.150000 ;
        RECT 1158.000000 287.850000 1168.000000 288.150000 ;
        RECT 1158.000000 291.850000 1168.000000 292.150000 ;
        RECT 1158.000000 295.850000 1168.000000 296.150000 ;
        RECT 1158.000000 299.850000 1168.000000 300.150000 ;
        RECT 1158.000000 303.850000 1168.000000 304.150000 ;
        RECT 1158.000000 307.850000 1168.000000 308.150000 ;
        RECT 1158.000000 311.850000 1168.000000 312.150000 ;
        RECT 1158.000000 315.850000 1168.000000 316.150000 ;
        RECT 1158.000000 319.850000 1168.000000 320.150000 ;
        RECT 1158.000000 323.850000 1168.000000 324.150000 ;
        RECT 1158.000000 339.850000 1168.000000 340.150000 ;
        RECT 1158.000000 335.850000 1168.000000 336.150000 ;
        RECT 1158.000000 331.850000 1168.000000 332.150000 ;
        RECT 1158.000000 327.850000 1168.000000 328.150000 ;
        RECT 60.000000 379.850000 65.000000 380.150000 ;
        RECT 18.000000 379.850000 28.000000 380.150000 ;
        RECT 18.000000 343.850000 28.000000 344.150000 ;
        RECT 18.000000 347.850000 28.000000 348.150000 ;
        RECT 18.000000 351.850000 28.000000 352.150000 ;
        RECT 18.000000 359.850000 28.000000 360.150000 ;
        RECT 18.000000 355.850000 28.000000 356.150000 ;
        RECT 18.000000 375.850000 28.000000 376.150000 ;
        RECT 18.000000 371.850000 28.000000 372.150000 ;
        RECT 18.000000 367.850000 28.000000 368.150000 ;
        RECT 18.000000 363.850000 28.000000 364.150000 ;
        RECT 60.000000 347.850000 65.000000 348.150000 ;
        RECT 60.000000 343.850000 65.000000 344.150000 ;
        RECT 60.000000 352.445000 64.080000 352.745000 ;
        RECT 60.000000 375.850000 65.000000 376.150000 ;
        RECT 60.000000 371.850000 65.000000 372.150000 ;
        RECT 60.000000 367.850000 65.000000 368.150000 ;
        RECT 60.000000 363.850000 65.000000 364.150000 ;
        RECT 18.000000 395.850000 28.000000 396.150000 ;
        RECT 18.000000 391.850000 28.000000 392.150000 ;
        RECT 18.000000 387.850000 28.000000 388.150000 ;
        RECT 18.000000 383.850000 28.000000 384.150000 ;
        RECT 18.000000 407.850000 28.000000 408.150000 ;
        RECT 18.000000 399.850000 28.000000 400.150000 ;
        RECT 18.000000 403.850000 28.000000 404.150000 ;
        RECT 18.000000 411.850000 28.000000 412.150000 ;
        RECT 18.000000 415.850000 28.000000 416.150000 ;
        RECT 60.000000 395.850000 65.000000 396.150000 ;
        RECT 60.000000 391.850000 65.000000 392.150000 ;
        RECT 60.000000 387.850000 65.000000 388.150000 ;
        RECT 60.000000 383.850000 65.000000 384.150000 ;
        RECT 60.000000 407.850000 65.000000 408.150000 ;
        RECT 60.000000 399.850000 65.000000 400.150000 ;
        RECT 60.000000 403.850000 65.000000 404.150000 ;
        RECT 60.000000 411.850000 65.000000 412.150000 ;
        RECT 60.000000 415.850000 65.000000 416.150000 ;
        RECT 110.000000 379.850000 115.000000 380.150000 ;
        RECT 110.000000 351.850000 115.000000 352.150000 ;
        RECT 110.000000 347.850000 115.000000 348.150000 ;
        RECT 110.000000 343.850000 115.000000 344.150000 ;
        RECT 110.000000 359.850000 115.000000 360.150000 ;
        RECT 110.000000 355.850000 115.000000 356.150000 ;
        RECT 110.000000 375.850000 115.000000 376.150000 ;
        RECT 110.000000 371.850000 115.000000 372.150000 ;
        RECT 110.000000 367.850000 115.000000 368.150000 ;
        RECT 110.000000 363.850000 115.000000 364.150000 ;
        RECT 110.000000 383.850000 115.000000 384.150000 ;
        RECT 110.000000 387.850000 115.000000 388.150000 ;
        RECT 110.000000 391.850000 115.000000 392.150000 ;
        RECT 110.000000 395.850000 115.000000 396.150000 ;
        RECT 110.000000 407.850000 115.000000 408.150000 ;
        RECT 110.000000 399.850000 115.000000 400.150000 ;
        RECT 110.000000 403.850000 115.000000 404.150000 ;
        RECT 110.000000 411.850000 115.000000 412.150000 ;
        RECT 110.000000 415.850000 115.000000 416.150000 ;
        RECT 18.000000 431.850000 28.000000 432.150000 ;
        RECT 18.000000 427.850000 28.000000 428.150000 ;
        RECT 18.000000 423.850000 28.000000 424.150000 ;
        RECT 18.000000 419.850000 28.000000 420.150000 ;
        RECT 18.000000 435.850000 28.000000 436.150000 ;
        RECT 18.000000 439.850000 28.000000 440.150000 ;
        RECT 18.000000 443.850000 28.000000 444.150000 ;
        RECT 18.000000 447.850000 28.000000 448.150000 ;
        RECT 18.000000 451.850000 28.000000 452.150000 ;
        RECT 60.000000 431.850000 65.000000 432.150000 ;
        RECT 60.000000 427.850000 65.000000 428.150000 ;
        RECT 60.000000 423.850000 65.000000 424.150000 ;
        RECT 60.000000 419.850000 65.000000 420.150000 ;
        RECT 60.000000 435.850000 65.000000 436.150000 ;
        RECT 60.000000 439.850000 65.000000 440.150000 ;
        RECT 60.000000 443.850000 65.000000 444.150000 ;
        RECT 60.000000 447.850000 65.000000 448.150000 ;
        RECT 60.000000 451.850000 65.000000 452.150000 ;
        RECT 18.000000 455.850000 28.000000 456.150000 ;
        RECT 18.000000 459.850000 28.000000 460.150000 ;
        RECT 18.000000 463.850000 28.000000 464.150000 ;
        RECT 18.000000 467.850000 28.000000 468.150000 ;
        RECT 18.000000 471.850000 28.000000 472.150000 ;
        RECT 18.000000 487.850000 28.000000 488.150000 ;
        RECT 18.000000 483.850000 28.000000 484.150000 ;
        RECT 18.000000 479.850000 28.000000 480.150000 ;
        RECT 18.000000 475.850000 28.000000 476.150000 ;
        RECT 60.000000 455.850000 65.000000 456.150000 ;
        RECT 60.000000 459.850000 65.000000 460.150000 ;
        RECT 60.000000 463.850000 65.000000 464.150000 ;
        RECT 60.000000 467.850000 65.000000 468.150000 ;
        RECT 60.000000 471.850000 65.000000 472.150000 ;
        RECT 60.000000 487.850000 65.000000 488.150000 ;
        RECT 60.000000 483.850000 65.000000 484.150000 ;
        RECT 60.000000 479.850000 65.000000 480.150000 ;
        RECT 60.000000 475.850000 65.000000 476.150000 ;
        RECT 110.000000 419.850000 115.000000 420.150000 ;
        RECT 110.000000 423.850000 115.000000 424.150000 ;
        RECT 110.000000 427.850000 115.000000 428.150000 ;
        RECT 110.000000 431.850000 115.000000 432.150000 ;
        RECT 110.000000 435.850000 115.000000 436.150000 ;
        RECT 110.000000 439.850000 115.000000 440.150000 ;
        RECT 110.000000 443.850000 115.000000 444.150000 ;
        RECT 110.000000 447.850000 115.000000 448.150000 ;
        RECT 110.000000 451.850000 115.000000 452.150000 ;
        RECT 110.000000 459.850000 115.000000 460.150000 ;
        RECT 110.000000 455.850000 115.000000 456.150000 ;
        RECT 110.000000 471.850000 115.000000 472.150000 ;
        RECT 110.000000 467.850000 115.000000 468.150000 ;
        RECT 110.000000 463.850000 115.000000 464.150000 ;
        RECT 110.000000 487.850000 115.000000 488.150000 ;
        RECT 110.000000 483.850000 115.000000 484.150000 ;
        RECT 110.000000 479.850000 115.000000 480.150000 ;
        RECT 110.000000 475.850000 115.000000 476.150000 ;
        RECT 210.000000 379.850000 215.000000 380.150000 ;
        RECT 160.000000 379.850000 165.000000 380.150000 ;
        RECT 160.000000 343.850000 165.000000 344.150000 ;
        RECT 160.000000 347.850000 165.000000 348.150000 ;
        RECT 160.000000 351.850000 165.000000 352.150000 ;
        RECT 160.000000 359.850000 165.000000 360.150000 ;
        RECT 160.000000 355.850000 165.000000 356.150000 ;
        RECT 160.000000 363.850000 165.000000 364.150000 ;
        RECT 160.000000 367.850000 165.000000 368.150000 ;
        RECT 160.000000 371.850000 165.000000 372.150000 ;
        RECT 160.000000 375.850000 165.000000 376.150000 ;
        RECT 210.000000 343.850000 215.000000 344.150000 ;
        RECT 210.000000 347.850000 215.000000 348.150000 ;
        RECT 210.000000 351.850000 215.000000 352.150000 ;
        RECT 210.000000 355.850000 215.000000 356.150000 ;
        RECT 210.000000 359.850000 215.000000 360.150000 ;
        RECT 210.000000 375.850000 215.000000 376.150000 ;
        RECT 210.000000 371.850000 215.000000 372.150000 ;
        RECT 210.000000 367.850000 215.000000 368.150000 ;
        RECT 210.000000 363.850000 215.000000 364.150000 ;
        RECT 160.000000 387.850000 165.000000 388.150000 ;
        RECT 160.000000 383.850000 165.000000 384.150000 ;
        RECT 160.000000 391.850000 165.000000 392.150000 ;
        RECT 160.000000 395.850000 165.000000 396.150000 ;
        RECT 160.000000 399.850000 165.000000 400.150000 ;
        RECT 210.000000 383.850000 215.000000 384.150000 ;
        RECT 210.000000 387.850000 215.000000 388.150000 ;
        RECT 210.000000 391.850000 215.000000 392.150000 ;
        RECT 210.000000 395.850000 215.000000 396.150000 ;
        RECT 210.000000 407.850000 215.000000 408.150000 ;
        RECT 210.000000 399.850000 215.000000 400.150000 ;
        RECT 210.000000 403.850000 215.000000 404.150000 ;
        RECT 210.000000 411.850000 215.000000 412.150000 ;
        RECT 210.000000 415.850000 215.000000 416.150000 ;
        RECT 260.000000 379.850000 265.000000 380.150000 ;
        RECT 260.000000 343.850000 265.000000 344.150000 ;
        RECT 260.000000 347.850000 265.000000 348.150000 ;
        RECT 260.000000 351.850000 265.000000 352.150000 ;
        RECT 260.000000 355.850000 265.000000 356.150000 ;
        RECT 260.000000 359.850000 265.000000 360.150000 ;
        RECT 260.000000 363.850000 265.000000 364.150000 ;
        RECT 260.000000 367.850000 265.000000 368.150000 ;
        RECT 260.000000 371.850000 265.000000 372.150000 ;
        RECT 260.000000 375.850000 265.000000 376.150000 ;
        RECT 260.000000 383.850000 265.000000 384.150000 ;
        RECT 260.000000 387.850000 265.000000 388.150000 ;
        RECT 260.000000 391.850000 265.000000 392.150000 ;
        RECT 260.000000 395.850000 265.000000 396.150000 ;
        RECT 260.000000 399.850000 265.000000 400.150000 ;
        RECT 210.000000 431.850000 215.000000 432.150000 ;
        RECT 210.000000 427.850000 215.000000 428.150000 ;
        RECT 210.000000 423.850000 215.000000 424.150000 ;
        RECT 210.000000 419.850000 215.000000 420.150000 ;
        RECT 210.000000 435.850000 215.000000 436.150000 ;
        RECT 210.000000 439.850000 215.000000 440.150000 ;
        RECT 210.000000 443.850000 215.000000 444.150000 ;
        RECT 210.000000 447.850000 215.000000 448.150000 ;
        RECT 210.000000 451.850000 215.000000 452.150000 ;
        RECT 160.000000 463.850000 165.000000 464.150000 ;
        RECT 160.000000 467.850000 165.000000 468.150000 ;
        RECT 160.000000 471.850000 165.000000 472.150000 ;
        RECT 160.000000 479.850000 165.000000 480.150000 ;
        RECT 160.000000 475.850000 165.000000 476.150000 ;
        RECT 160.000000 487.850000 165.000000 488.150000 ;
        RECT 160.000000 483.850000 165.000000 484.150000 ;
        RECT 210.000000 455.850000 215.000000 456.150000 ;
        RECT 210.000000 459.850000 215.000000 460.150000 ;
        RECT 210.000000 463.850000 215.000000 464.150000 ;
        RECT 210.000000 467.850000 215.000000 468.150000 ;
        RECT 210.000000 471.850000 215.000000 472.150000 ;
        RECT 210.000000 475.850000 215.000000 476.150000 ;
        RECT 210.000000 479.850000 215.000000 480.150000 ;
        RECT 210.000000 483.850000 215.000000 484.150000 ;
        RECT 210.000000 487.850000 215.000000 488.150000 ;
        RECT 260.000000 467.850000 265.000000 468.150000 ;
        RECT 260.000000 463.850000 265.000000 464.150000 ;
        RECT 260.000000 471.850000 265.000000 472.150000 ;
        RECT 260.000000 475.850000 265.000000 476.150000 ;
        RECT 260.000000 479.850000 265.000000 480.150000 ;
        RECT 260.000000 487.850000 265.000000 488.150000 ;
        RECT 260.000000 483.850000 265.000000 484.150000 ;
        RECT 18.000000 491.850000 28.000000 492.150000 ;
        RECT 18.000000 495.850000 28.000000 496.150000 ;
        RECT 18.000000 499.850000 28.000000 500.150000 ;
        RECT 18.000000 503.850000 28.000000 504.150000 ;
        RECT 18.000000 507.850000 28.000000 508.150000 ;
        RECT 18.000000 515.850000 28.000000 516.150000 ;
        RECT 18.000000 511.850000 28.000000 512.150000 ;
        RECT 60.000000 491.850000 65.000000 492.150000 ;
        RECT 60.000000 495.850000 65.000000 496.150000 ;
        RECT 60.000000 499.850000 65.000000 500.150000 ;
        RECT 60.000000 503.850000 65.000000 504.150000 ;
        RECT 60.000000 507.850000 65.000000 508.150000 ;
        RECT 60.000000 515.850000 65.000000 516.150000 ;
        RECT 60.000000 511.850000 65.000000 512.150000 ;
        RECT 110.000000 499.850000 115.000000 500.150000 ;
        RECT 110.000000 495.850000 115.000000 496.150000 ;
        RECT 110.000000 491.850000 115.000000 492.150000 ;
        RECT 110.000000 507.850000 115.000000 508.150000 ;
        RECT 110.000000 503.850000 115.000000 504.150000 ;
        RECT 110.000000 515.850000 115.000000 516.150000 ;
        RECT 110.000000 511.850000 115.000000 512.150000 ;
        RECT 160.000000 491.850000 165.000000 492.150000 ;
        RECT 160.000000 495.850000 165.000000 496.150000 ;
        RECT 160.000000 499.850000 165.000000 500.150000 ;
        RECT 160.000000 507.850000 165.000000 508.150000 ;
        RECT 160.000000 503.850000 165.000000 504.150000 ;
        RECT 160.000000 515.850000 165.000000 516.150000 ;
        RECT 160.000000 511.850000 165.000000 512.150000 ;
        RECT 210.000000 491.850000 215.000000 492.150000 ;
        RECT 210.000000 495.850000 215.000000 496.150000 ;
        RECT 210.000000 499.850000 215.000000 500.150000 ;
        RECT 210.000000 503.850000 215.000000 504.150000 ;
        RECT 210.000000 507.850000 215.000000 508.150000 ;
        RECT 210.000000 515.850000 215.000000 516.150000 ;
        RECT 210.000000 511.850000 215.000000 512.150000 ;
        RECT 260.000000 495.850000 265.000000 496.150000 ;
        RECT 260.000000 491.850000 265.000000 492.150000 ;
        RECT 260.000000 499.850000 265.000000 500.150000 ;
        RECT 260.000000 507.850000 265.000000 508.150000 ;
        RECT 260.000000 503.850000 265.000000 504.150000 ;
        RECT 260.000000 515.850000 265.000000 516.150000 ;
        RECT 260.000000 511.850000 265.000000 512.150000 ;
        RECT 360.000000 379.850000 365.000000 380.150000 ;
        RECT 310.000000 379.850000 315.000000 380.150000 ;
        RECT 310.000000 343.850000 315.000000 344.150000 ;
        RECT 310.000000 351.850000 315.000000 352.150000 ;
        RECT 310.000000 347.850000 315.000000 348.150000 ;
        RECT 310.000000 355.850000 315.000000 356.150000 ;
        RECT 310.000000 359.850000 315.000000 360.150000 ;
        RECT 310.000000 363.850000 315.000000 364.150000 ;
        RECT 310.000000 367.850000 315.000000 368.150000 ;
        RECT 310.000000 371.850000 315.000000 372.150000 ;
        RECT 310.000000 375.850000 315.000000 376.150000 ;
        RECT 360.000000 343.850000 365.000000 344.150000 ;
        RECT 360.000000 347.850000 365.000000 348.150000 ;
        RECT 360.000000 351.850000 365.000000 352.150000 ;
        RECT 360.000000 355.850000 365.000000 356.150000 ;
        RECT 360.000000 359.850000 365.000000 360.150000 ;
        RECT 360.000000 375.850000 365.000000 376.150000 ;
        RECT 360.000000 371.850000 365.000000 372.150000 ;
        RECT 360.000000 367.850000 365.000000 368.150000 ;
        RECT 360.000000 363.850000 365.000000 364.150000 ;
        RECT 310.000000 383.850000 315.000000 384.150000 ;
        RECT 310.000000 387.850000 315.000000 388.150000 ;
        RECT 310.000000 391.850000 315.000000 392.150000 ;
        RECT 310.000000 395.850000 315.000000 396.150000 ;
        RECT 310.000000 407.850000 315.000000 408.150000 ;
        RECT 310.000000 399.850000 315.000000 400.150000 ;
        RECT 310.000000 403.850000 315.000000 404.150000 ;
        RECT 310.000000 411.850000 315.000000 412.150000 ;
        RECT 310.000000 415.850000 315.000000 416.150000 ;
        RECT 360.000000 383.850000 365.000000 384.150000 ;
        RECT 360.000000 387.850000 365.000000 388.150000 ;
        RECT 360.000000 391.850000 365.000000 392.150000 ;
        RECT 360.000000 395.850000 365.000000 396.150000 ;
        RECT 360.000000 407.850000 365.000000 408.150000 ;
        RECT 360.000000 399.850000 365.000000 400.150000 ;
        RECT 360.000000 403.850000 365.000000 404.150000 ;
        RECT 360.000000 411.850000 365.000000 412.150000 ;
        RECT 360.000000 415.850000 365.000000 416.150000 ;
        RECT 410.000000 379.850000 415.000000 380.150000 ;
        RECT 410.000000 351.850000 415.000000 352.150000 ;
        RECT 410.000000 347.850000 415.000000 348.150000 ;
        RECT 410.000000 343.850000 415.000000 344.150000 ;
        RECT 410.000000 355.850000 415.000000 356.150000 ;
        RECT 410.000000 359.850000 415.000000 360.150000 ;
        RECT 410.000000 375.850000 415.000000 376.150000 ;
        RECT 410.000000 371.850000 415.000000 372.150000 ;
        RECT 410.000000 367.850000 415.000000 368.150000 ;
        RECT 410.000000 363.850000 415.000000 364.150000 ;
        RECT 410.000000 383.850000 415.000000 384.150000 ;
        RECT 410.000000 387.850000 415.000000 388.150000 ;
        RECT 410.000000 391.850000 415.000000 392.150000 ;
        RECT 410.000000 395.850000 415.000000 396.150000 ;
        RECT 410.000000 407.850000 415.000000 408.150000 ;
        RECT 410.000000 399.850000 415.000000 400.150000 ;
        RECT 410.000000 403.850000 415.000000 404.150000 ;
        RECT 410.000000 411.850000 415.000000 412.150000 ;
        RECT 410.000000 415.850000 415.000000 416.150000 ;
        RECT 310.000000 419.850000 315.000000 420.150000 ;
        RECT 310.000000 423.850000 315.000000 424.150000 ;
        RECT 310.000000 427.850000 315.000000 428.150000 ;
        RECT 310.000000 431.850000 315.000000 432.150000 ;
        RECT 310.000000 439.850000 315.000000 440.150000 ;
        RECT 310.000000 435.850000 315.000000 436.150000 ;
        RECT 310.000000 443.850000 315.000000 444.150000 ;
        RECT 310.000000 447.850000 315.000000 448.150000 ;
        RECT 310.000000 451.850000 315.000000 452.150000 ;
        RECT 360.000000 419.850000 365.000000 420.150000 ;
        RECT 360.000000 423.850000 365.000000 424.150000 ;
        RECT 360.000000 427.850000 365.000000 428.150000 ;
        RECT 360.000000 431.850000 365.000000 432.150000 ;
        RECT 360.000000 435.850000 365.000000 436.150000 ;
        RECT 360.000000 439.850000 365.000000 440.150000 ;
        RECT 360.000000 443.850000 365.000000 444.150000 ;
        RECT 360.000000 447.850000 365.000000 448.150000 ;
        RECT 360.000000 451.850000 365.000000 452.150000 ;
        RECT 310.000000 459.850000 315.000000 460.150000 ;
        RECT 310.000000 455.850000 315.000000 456.150000 ;
        RECT 310.000000 467.850000 315.000000 468.150000 ;
        RECT 310.000000 463.850000 315.000000 464.150000 ;
        RECT 310.000000 471.850000 315.000000 472.150000 ;
        RECT 310.000000 475.850000 315.000000 476.150000 ;
        RECT 310.000000 479.850000 315.000000 480.150000 ;
        RECT 310.000000 483.850000 315.000000 484.150000 ;
        RECT 310.000000 487.850000 315.000000 488.150000 ;
        RECT 360.000000 455.850000 365.000000 456.150000 ;
        RECT 360.000000 459.850000 365.000000 460.150000 ;
        RECT 360.000000 463.850000 365.000000 464.150000 ;
        RECT 360.000000 467.850000 365.000000 468.150000 ;
        RECT 360.000000 471.850000 365.000000 472.150000 ;
        RECT 360.000000 475.850000 365.000000 476.150000 ;
        RECT 360.000000 479.850000 365.000000 480.150000 ;
        RECT 360.000000 483.850000 365.000000 484.150000 ;
        RECT 360.000000 487.850000 365.000000 488.150000 ;
        RECT 410.000000 423.850000 415.000000 424.150000 ;
        RECT 410.000000 419.850000 415.000000 420.150000 ;
        RECT 410.000000 427.850000 415.000000 428.150000 ;
        RECT 410.000000 431.850000 415.000000 432.150000 ;
        RECT 410.000000 439.850000 415.000000 440.150000 ;
        RECT 410.000000 435.850000 415.000000 436.150000 ;
        RECT 410.000000 443.850000 415.000000 444.150000 ;
        RECT 410.000000 447.850000 415.000000 448.150000 ;
        RECT 410.000000 451.850000 415.000000 452.150000 ;
        RECT 371.000000 479.850000 381.000000 480.150000 ;
        RECT 371.000000 483.850000 381.000000 484.150000 ;
        RECT 371.000000 487.850000 381.000000 488.150000 ;
        RECT 410.000000 455.850000 415.000000 456.150000 ;
        RECT 410.000000 459.850000 415.000000 460.150000 ;
        RECT 410.000000 467.850000 415.000000 468.150000 ;
        RECT 410.000000 463.850000 415.000000 464.150000 ;
        RECT 410.000000 471.850000 415.000000 472.150000 ;
        RECT 410.000000 475.850000 415.000000 476.150000 ;
        RECT 410.000000 479.850000 415.000000 480.150000 ;
        RECT 410.000000 483.850000 415.000000 484.150000 ;
        RECT 410.000000 487.850000 415.000000 488.150000 ;
        RECT 460.000000 379.850000 465.000000 380.150000 ;
        RECT 510.000000 379.850000 515.000000 380.150000 ;
        RECT 460.000000 347.850000 465.000000 348.150000 ;
        RECT 460.000000 343.850000 465.000000 344.150000 ;
        RECT 460.000000 351.230000 465.000000 352.230000 ;
        RECT 460.000000 375.850000 465.000000 376.150000 ;
        RECT 460.000000 371.850000 465.000000 372.150000 ;
        RECT 510.000000 343.850000 515.000000 344.150000 ;
        RECT 510.000000 351.850000 515.000000 352.150000 ;
        RECT 510.000000 347.850000 515.000000 348.150000 ;
        RECT 510.000000 359.850000 515.000000 360.150000 ;
        RECT 510.000000 355.850000 515.000000 356.150000 ;
        RECT 510.000000 363.850000 515.000000 364.150000 ;
        RECT 510.000000 367.850000 515.000000 368.150000 ;
        RECT 510.000000 375.850000 515.000000 376.150000 ;
        RECT 510.000000 371.850000 515.000000 372.150000 ;
        RECT 460.000000 395.850000 465.000000 396.150000 ;
        RECT 460.000000 391.850000 465.000000 392.150000 ;
        RECT 460.000000 387.850000 465.000000 388.150000 ;
        RECT 460.000000 383.850000 465.000000 384.150000 ;
        RECT 460.000000 401.230000 465.000000 402.230000 ;
        RECT 510.000000 383.850000 515.000000 384.150000 ;
        RECT 510.000000 387.850000 515.000000 388.150000 ;
        RECT 510.000000 391.850000 515.000000 392.150000 ;
        RECT 510.000000 395.850000 515.000000 396.150000 ;
        RECT 510.000000 407.850000 515.000000 408.150000 ;
        RECT 510.000000 399.850000 515.000000 400.150000 ;
        RECT 510.000000 403.850000 515.000000 404.150000 ;
        RECT 510.000000 411.850000 515.000000 412.150000 ;
        RECT 510.000000 415.850000 515.000000 416.150000 ;
        RECT 560.000000 379.850000 565.000000 380.150000 ;
        RECT 560.000000 359.850000 565.000000 360.150000 ;
        RECT 560.000000 355.850000 565.000000 356.150000 ;
        RECT 560.000000 351.850000 565.000000 352.150000 ;
        RECT 560.000000 347.850000 565.000000 348.150000 ;
        RECT 560.000000 343.850000 565.000000 344.150000 ;
        RECT 560.000000 375.850000 565.000000 376.150000 ;
        RECT 560.000000 371.850000 565.000000 372.150000 ;
        RECT 560.000000 367.850000 565.000000 368.150000 ;
        RECT 560.000000 363.850000 565.000000 364.150000 ;
        RECT 560.000000 383.850000 565.000000 384.150000 ;
        RECT 560.000000 387.850000 565.000000 388.150000 ;
        RECT 560.000000 395.850000 565.000000 396.150000 ;
        RECT 560.000000 391.850000 565.000000 392.150000 ;
        RECT 560.000000 407.850000 565.000000 408.150000 ;
        RECT 560.000000 399.850000 565.000000 400.150000 ;
        RECT 560.000000 403.850000 565.000000 404.150000 ;
        RECT 560.000000 415.850000 565.000000 416.150000 ;
        RECT 560.000000 411.850000 565.000000 412.150000 ;
        RECT 460.000000 419.850000 465.000000 420.150000 ;
        RECT 460.000000 423.850000 465.000000 424.150000 ;
        RECT 460.000000 427.850000 465.000000 428.150000 ;
        RECT 460.000000 431.850000 465.000000 432.150000 ;
        RECT 460.000000 435.850000 465.000000 436.150000 ;
        RECT 460.000000 439.850000 465.000000 440.150000 ;
        RECT 460.000000 443.850000 465.000000 444.150000 ;
        RECT 460.000000 447.850000 465.000000 448.150000 ;
        RECT 460.000000 451.850000 465.000000 452.150000 ;
        RECT 510.000000 419.850000 515.000000 420.150000 ;
        RECT 510.000000 423.850000 515.000000 424.150000 ;
        RECT 510.000000 427.850000 515.000000 428.150000 ;
        RECT 510.000000 431.850000 515.000000 432.150000 ;
        RECT 510.000000 439.850000 515.000000 440.150000 ;
        RECT 510.000000 435.850000 515.000000 436.150000 ;
        RECT 510.000000 443.850000 515.000000 444.150000 ;
        RECT 510.000000 447.850000 515.000000 448.150000 ;
        RECT 510.000000 451.850000 515.000000 452.150000 ;
        RECT 460.000000 455.850000 465.000000 456.150000 ;
        RECT 460.000000 459.850000 465.000000 460.150000 ;
        RECT 460.000000 463.850000 465.000000 464.150000 ;
        RECT 460.000000 467.850000 465.000000 468.150000 ;
        RECT 460.000000 471.850000 465.000000 472.150000 ;
        RECT 460.000000 475.850000 465.000000 476.150000 ;
        RECT 460.000000 479.850000 465.000000 480.150000 ;
        RECT 460.000000 483.850000 465.000000 484.150000 ;
        RECT 460.000000 487.850000 465.000000 488.150000 ;
        RECT 510.000000 455.850000 515.000000 456.150000 ;
        RECT 510.000000 459.850000 515.000000 460.150000 ;
        RECT 510.000000 467.850000 515.000000 468.150000 ;
        RECT 510.000000 463.850000 515.000000 464.150000 ;
        RECT 510.000000 471.850000 515.000000 472.150000 ;
        RECT 510.000000 475.850000 515.000000 476.150000 ;
        RECT 510.000000 479.850000 515.000000 480.150000 ;
        RECT 510.000000 483.850000 515.000000 484.150000 ;
        RECT 510.000000 487.850000 515.000000 488.150000 ;
        RECT 560.000000 423.850000 565.000000 424.150000 ;
        RECT 560.000000 419.850000 565.000000 420.150000 ;
        RECT 560.000000 427.850000 565.000000 428.150000 ;
        RECT 560.000000 431.850000 565.000000 432.150000 ;
        RECT 560.000000 435.850000 565.000000 436.150000 ;
        RECT 560.000000 439.850000 565.000000 440.150000 ;
        RECT 560.000000 443.850000 565.000000 444.150000 ;
        RECT 560.000000 447.850000 565.000000 448.150000 ;
        RECT 560.000000 451.850000 565.000000 452.150000 ;
        RECT 560.000000 455.850000 565.000000 456.150000 ;
        RECT 560.000000 459.850000 565.000000 460.150000 ;
        RECT 560.000000 467.850000 565.000000 468.150000 ;
        RECT 560.000000 463.850000 565.000000 464.150000 ;
        RECT 560.000000 471.850000 565.000000 472.150000 ;
        RECT 560.000000 475.850000 565.000000 476.150000 ;
        RECT 560.000000 479.850000 565.000000 480.150000 ;
        RECT 560.000000 483.850000 565.000000 484.150000 ;
        RECT 560.000000 487.850000 565.000000 488.150000 ;
        RECT 310.000000 495.850000 315.000000 496.150000 ;
        RECT 310.000000 491.850000 315.000000 492.150000 ;
        RECT 310.000000 499.850000 315.000000 500.150000 ;
        RECT 310.000000 507.850000 315.000000 508.150000 ;
        RECT 310.000000 503.850000 315.000000 504.150000 ;
        RECT 310.000000 515.850000 315.000000 516.150000 ;
        RECT 310.000000 511.850000 315.000000 512.150000 ;
        RECT 360.000000 491.850000 365.000000 492.150000 ;
        RECT 360.000000 495.850000 365.000000 496.150000 ;
        RECT 360.000000 499.850000 365.000000 500.150000 ;
        RECT 360.000000 503.850000 365.000000 504.150000 ;
        RECT 360.000000 507.850000 365.000000 508.150000 ;
        RECT 360.000000 511.850000 365.000000 512.150000 ;
        RECT 360.000000 515.850000 365.000000 516.150000 ;
        RECT 360.000000 519.850000 365.000000 520.150000 ;
        RECT 360.000000 523.850000 365.000000 524.150000 ;
        RECT 360.000000 527.850000 365.000000 528.150000 ;
        RECT 360.000000 531.850000 365.000000 532.150000 ;
        RECT 360.000000 535.850000 365.000000 536.150000 ;
        RECT 360.000000 539.850000 365.000000 540.150000 ;
        RECT 360.000000 543.850000 365.000000 544.150000 ;
        RECT 360.000000 555.850000 365.000000 556.150000 ;
        RECT 360.000000 547.850000 365.000000 548.150000 ;
        RECT 360.000000 551.850000 365.000000 552.150000 ;
        RECT 360.000000 559.850000 365.000000 560.150000 ;
        RECT 360.000000 563.850000 365.000000 564.150000 ;
        RECT 371.000000 491.850000 381.000000 492.150000 ;
        RECT 371.000000 495.850000 381.000000 496.150000 ;
        RECT 371.000000 499.850000 381.000000 500.150000 ;
        RECT 371.000000 503.850000 381.000000 504.150000 ;
        RECT 371.000000 507.850000 381.000000 508.150000 ;
        RECT 371.000000 511.850000 381.000000 512.150000 ;
        RECT 371.000000 515.850000 381.000000 516.150000 ;
        RECT 371.000000 519.850000 381.000000 520.150000 ;
        RECT 371.000000 523.850000 381.000000 524.150000 ;
        RECT 371.000000 527.850000 381.000000 528.150000 ;
        RECT 410.000000 495.850000 415.000000 496.150000 ;
        RECT 410.000000 491.850000 415.000000 492.150000 ;
        RECT 410.000000 499.850000 415.000000 500.150000 ;
        RECT 410.000000 503.850000 415.000000 504.150000 ;
        RECT 371.000000 531.850000 381.000000 532.150000 ;
        RECT 371.000000 535.850000 381.000000 536.150000 ;
        RECT 371.000000 539.850000 381.000000 540.150000 ;
        RECT 371.000000 543.850000 381.000000 544.150000 ;
        RECT 371.000000 555.850000 381.000000 556.150000 ;
        RECT 371.000000 547.850000 381.000000 548.150000 ;
        RECT 371.000000 551.850000 381.000000 552.150000 ;
        RECT 371.000000 559.850000 381.000000 560.150000 ;
        RECT 371.000000 563.850000 381.000000 564.150000 ;
        RECT 360.000000 583.850000 365.000000 584.150000 ;
        RECT 360.000000 567.850000 365.000000 568.150000 ;
        RECT 360.000000 571.850000 365.000000 572.150000 ;
        RECT 360.000000 575.850000 365.000000 576.150000 ;
        RECT 360.000000 579.850000 365.000000 580.150000 ;
        RECT 360.000000 587.850000 365.000000 588.150000 ;
        RECT 360.000000 591.850000 365.000000 592.150000 ;
        RECT 360.000000 595.850000 365.000000 596.150000 ;
        RECT 360.000000 599.850000 365.000000 600.150000 ;
        RECT 360.000000 603.850000 365.000000 604.150000 ;
        RECT 360.000000 607.850000 365.000000 608.150000 ;
        RECT 360.000000 611.850000 365.000000 612.150000 ;
        RECT 360.000000 615.850000 365.000000 616.150000 ;
        RECT 360.000000 619.850000 365.000000 620.150000 ;
        RECT 360.000000 623.850000 365.000000 624.150000 ;
        RECT 360.000000 627.850000 365.000000 628.150000 ;
        RECT 360.000000 631.850000 365.000000 632.150000 ;
        RECT 360.000000 635.850000 365.000000 636.150000 ;
        RECT 371.000000 583.850000 381.000000 584.150000 ;
        RECT 371.000000 579.850000 381.000000 580.150000 ;
        RECT 371.000000 575.850000 381.000000 576.150000 ;
        RECT 371.000000 571.850000 381.000000 572.150000 ;
        RECT 371.000000 567.850000 381.000000 568.150000 ;
        RECT 371.000000 587.850000 381.000000 588.150000 ;
        RECT 371.000000 591.850000 381.000000 592.150000 ;
        RECT 371.000000 595.850000 381.000000 596.150000 ;
        RECT 371.000000 599.850000 381.000000 600.150000 ;
        RECT 371.000000 603.850000 381.000000 604.150000 ;
        RECT 371.000000 607.850000 381.000000 608.150000 ;
        RECT 371.000000 611.850000 381.000000 612.150000 ;
        RECT 371.000000 615.850000 381.000000 616.150000 ;
        RECT 371.000000 619.850000 381.000000 620.150000 ;
        RECT 371.000000 635.850000 381.000000 636.150000 ;
        RECT 371.000000 631.850000 381.000000 632.150000 ;
        RECT 371.000000 627.850000 381.000000 628.150000 ;
        RECT 371.000000 623.850000 381.000000 624.150000 ;
        RECT 460.000000 495.850000 465.000000 496.150000 ;
        RECT 460.000000 491.850000 465.000000 492.150000 ;
        RECT 460.000000 499.850000 465.000000 500.150000 ;
        RECT 460.000000 503.850000 465.000000 504.150000 ;
        RECT 510.000000 495.850000 515.000000 496.150000 ;
        RECT 510.000000 491.850000 515.000000 492.150000 ;
        RECT 510.000000 499.850000 515.000000 500.150000 ;
        RECT 510.000000 503.850000 515.000000 504.150000 ;
        RECT 560.000000 503.850000 565.000000 504.150000 ;
        RECT 560.000000 499.850000 565.000000 500.150000 ;
        RECT 560.000000 495.850000 565.000000 496.150000 ;
        RECT 560.000000 491.850000 565.000000 492.150000 ;
        RECT 360.000000 639.850000 365.000000 640.150000 ;
        RECT 360.000000 643.850000 365.000000 644.150000 ;
        RECT 360.000000 647.850000 365.000000 648.150000 ;
        RECT 360.000000 651.850000 365.000000 652.150000 ;
        RECT 360.000000 655.850000 365.000000 656.150000 ;
        RECT 360.000000 659.850000 365.000000 660.150000 ;
        RECT 360.000000 663.850000 365.000000 664.150000 ;
        RECT 360.000000 667.850000 365.000000 668.150000 ;
        RECT 360.000000 671.850000 365.000000 672.150000 ;
        RECT 360.000000 675.850000 365.000000 676.150000 ;
        RECT 310.000000 679.850000 315.000000 680.150000 ;
        RECT 310.000000 683.850000 315.000000 684.150000 ;
        RECT 360.000000 679.850000 365.000000 680.150000 ;
        RECT 360.000000 683.850000 365.000000 684.150000 ;
        RECT 371.000000 639.850000 381.000000 640.150000 ;
        RECT 371.000000 643.850000 381.000000 644.150000 ;
        RECT 371.000000 647.850000 381.000000 648.150000 ;
        RECT 371.000000 651.850000 381.000000 652.150000 ;
        RECT 371.000000 655.850000 381.000000 656.150000 ;
        RECT 371.000000 667.850000 381.000000 668.150000 ;
        RECT 371.000000 663.850000 381.000000 664.150000 ;
        RECT 371.000000 659.850000 381.000000 660.150000 ;
        RECT 410.000000 659.850000 415.000000 660.150000 ;
        RECT 410.000000 663.850000 415.000000 664.150000 ;
        RECT 410.000000 667.850000 415.000000 668.150000 ;
        RECT 410.000000 671.850000 415.000000 672.150000 ;
        RECT 410.000000 675.850000 415.000000 676.150000 ;
        RECT 410.000000 683.850000 415.000000 684.150000 ;
        RECT 410.000000 679.850000 415.000000 680.150000 ;
        RECT 460.000000 659.850000 465.000000 660.150000 ;
        RECT 460.000000 663.850000 465.000000 664.150000 ;
        RECT 460.000000 667.850000 465.000000 668.150000 ;
        RECT 460.000000 671.850000 465.000000 672.150000 ;
        RECT 460.000000 675.850000 465.000000 676.150000 ;
        RECT 510.000000 659.850000 515.000000 660.150000 ;
        RECT 510.000000 663.850000 515.000000 664.150000 ;
        RECT 510.000000 667.850000 515.000000 668.150000 ;
        RECT 510.000000 671.850000 515.000000 672.150000 ;
        RECT 510.000000 675.850000 515.000000 676.150000 ;
        RECT 460.000000 683.850000 465.000000 684.150000 ;
        RECT 460.000000 679.850000 465.000000 680.150000 ;
        RECT 510.000000 683.850000 515.000000 684.150000 ;
        RECT 510.000000 679.850000 515.000000 680.150000 ;
        RECT 560.000000 659.850000 565.000000 660.150000 ;
        RECT 560.000000 663.850000 565.000000 664.150000 ;
        RECT 560.000000 667.850000 565.000000 668.150000 ;
        RECT 560.000000 671.850000 565.000000 672.150000 ;
        RECT 560.000000 675.850000 565.000000 676.150000 ;
        RECT 560.000000 683.850000 565.000000 684.150000 ;
        RECT 560.000000 679.850000 565.000000 680.150000 ;
        RECT 610.000000 379.850000 615.000000 380.150000 ;
        RECT 660.000000 379.850000 665.000000 380.150000 ;
        RECT 610.000000 343.850000 615.000000 344.150000 ;
        RECT 610.000000 347.850000 615.000000 348.150000 ;
        RECT 610.000000 351.850000 615.000000 352.150000 ;
        RECT 610.000000 355.850000 615.000000 356.150000 ;
        RECT 610.000000 359.850000 615.000000 360.150000 ;
        RECT 610.000000 375.850000 615.000000 376.150000 ;
        RECT 610.000000 371.850000 615.000000 372.150000 ;
        RECT 610.000000 367.850000 615.000000 368.150000 ;
        RECT 610.000000 363.850000 615.000000 364.150000 ;
        RECT 660.000000 343.850000 665.000000 344.150000 ;
        RECT 660.000000 347.850000 665.000000 348.150000 ;
        RECT 660.000000 351.850000 665.000000 352.150000 ;
        RECT 660.000000 359.850000 665.000000 360.150000 ;
        RECT 660.000000 355.850000 665.000000 356.150000 ;
        RECT 660.000000 363.850000 665.000000 364.150000 ;
        RECT 660.000000 367.850000 665.000000 368.150000 ;
        RECT 660.000000 371.850000 665.000000 372.150000 ;
        RECT 660.000000 375.850000 665.000000 376.150000 ;
        RECT 610.000000 383.850000 615.000000 384.150000 ;
        RECT 610.000000 387.850000 615.000000 388.150000 ;
        RECT 610.000000 391.850000 615.000000 392.150000 ;
        RECT 610.000000 395.850000 615.000000 396.150000 ;
        RECT 610.000000 407.850000 615.000000 408.150000 ;
        RECT 610.000000 399.850000 615.000000 400.150000 ;
        RECT 610.000000 403.850000 615.000000 404.150000 ;
        RECT 610.000000 411.850000 615.000000 412.150000 ;
        RECT 610.000000 415.850000 615.000000 416.150000 ;
        RECT 660.000000 383.850000 665.000000 384.150000 ;
        RECT 660.000000 387.850000 665.000000 388.150000 ;
        RECT 660.000000 391.850000 665.000000 392.150000 ;
        RECT 660.000000 395.850000 665.000000 396.150000 ;
        RECT 660.000000 407.850000 665.000000 408.150000 ;
        RECT 660.000000 399.850000 665.000000 400.150000 ;
        RECT 660.000000 403.850000 665.000000 404.150000 ;
        RECT 660.000000 411.850000 665.000000 412.150000 ;
        RECT 660.000000 415.850000 665.000000 416.150000 ;
        RECT 710.000000 379.850000 715.000000 380.150000 ;
        RECT 710.000000 359.850000 715.000000 360.150000 ;
        RECT 710.000000 355.850000 715.000000 356.150000 ;
        RECT 710.000000 351.850000 715.000000 352.150000 ;
        RECT 710.000000 347.850000 715.000000 348.150000 ;
        RECT 710.000000 343.850000 715.000000 344.150000 ;
        RECT 710.000000 375.850000 715.000000 376.150000 ;
        RECT 710.000000 371.850000 715.000000 372.150000 ;
        RECT 710.000000 367.850000 715.000000 368.150000 ;
        RECT 710.000000 363.850000 715.000000 364.150000 ;
        RECT 710.000000 383.850000 715.000000 384.150000 ;
        RECT 710.000000 387.850000 715.000000 388.150000 ;
        RECT 710.000000 391.850000 715.000000 392.150000 ;
        RECT 710.000000 395.850000 715.000000 396.150000 ;
        RECT 710.000000 407.850000 715.000000 408.150000 ;
        RECT 710.000000 403.850000 715.000000 404.150000 ;
        RECT 710.000000 399.850000 715.000000 400.150000 ;
        RECT 710.000000 415.850000 715.000000 416.150000 ;
        RECT 710.000000 411.850000 715.000000 412.150000 ;
        RECT 610.000000 419.850000 615.000000 420.150000 ;
        RECT 610.000000 423.850000 615.000000 424.150000 ;
        RECT 610.000000 427.850000 615.000000 428.150000 ;
        RECT 610.000000 431.850000 615.000000 432.150000 ;
        RECT 610.000000 435.850000 615.000000 436.150000 ;
        RECT 610.000000 439.850000 615.000000 440.150000 ;
        RECT 610.000000 443.850000 615.000000 444.150000 ;
        RECT 610.000000 447.850000 615.000000 448.150000 ;
        RECT 610.000000 451.850000 615.000000 452.150000 ;
        RECT 660.000000 419.850000 665.000000 420.150000 ;
        RECT 660.000000 423.850000 665.000000 424.150000 ;
        RECT 660.000000 427.850000 665.000000 428.150000 ;
        RECT 660.000000 431.850000 665.000000 432.150000 ;
        RECT 660.000000 435.850000 665.000000 436.150000 ;
        RECT 660.000000 439.850000 665.000000 440.150000 ;
        RECT 660.000000 443.850000 665.000000 444.150000 ;
        RECT 660.000000 447.850000 665.000000 448.150000 ;
        RECT 660.000000 451.850000 665.000000 452.150000 ;
        RECT 610.000000 455.850000 615.000000 456.150000 ;
        RECT 610.000000 459.850000 615.000000 460.150000 ;
        RECT 610.000000 463.850000 615.000000 464.150000 ;
        RECT 610.000000 467.850000 615.000000 468.150000 ;
        RECT 610.000000 471.850000 615.000000 472.150000 ;
        RECT 610.000000 487.850000 615.000000 488.150000 ;
        RECT 610.000000 483.850000 615.000000 484.150000 ;
        RECT 610.000000 479.850000 615.000000 480.150000 ;
        RECT 610.000000 475.850000 615.000000 476.150000 ;
        RECT 660.000000 455.850000 665.000000 456.150000 ;
        RECT 660.000000 459.850000 665.000000 460.150000 ;
        RECT 660.000000 463.850000 665.000000 464.150000 ;
        RECT 660.000000 467.850000 665.000000 468.150000 ;
        RECT 660.000000 471.850000 665.000000 472.150000 ;
        RECT 660.000000 479.850000 665.000000 480.150000 ;
        RECT 660.000000 475.850000 665.000000 476.150000 ;
        RECT 660.000000 487.850000 665.000000 488.150000 ;
        RECT 660.000000 483.850000 665.000000 484.150000 ;
        RECT 721.000000 431.850000 731.000000 432.150000 ;
        RECT 721.000000 419.850000 731.000000 420.150000 ;
        RECT 721.000000 423.850000 731.000000 424.150000 ;
        RECT 721.000000 427.850000 731.000000 428.150000 ;
        RECT 710.000000 419.850000 715.000000 420.150000 ;
        RECT 710.000000 423.850000 715.000000 424.150000 ;
        RECT 710.000000 427.850000 715.000000 428.150000 ;
        RECT 710.000000 431.850000 715.000000 432.150000 ;
        RECT 721.000000 435.850000 731.000000 436.150000 ;
        RECT 721.000000 439.850000 731.000000 440.150000 ;
        RECT 721.000000 443.850000 731.000000 444.150000 ;
        RECT 721.000000 447.850000 731.000000 448.150000 ;
        RECT 721.000000 451.850000 731.000000 452.150000 ;
        RECT 710.000000 439.850000 715.000000 440.150000 ;
        RECT 710.000000 435.850000 715.000000 436.150000 ;
        RECT 710.000000 443.850000 715.000000 444.150000 ;
        RECT 710.000000 447.850000 715.000000 448.150000 ;
        RECT 710.000000 451.850000 715.000000 452.150000 ;
        RECT 721.000000 459.850000 731.000000 460.150000 ;
        RECT 721.000000 455.850000 731.000000 456.150000 ;
        RECT 721.000000 463.850000 731.000000 464.150000 ;
        RECT 721.000000 467.850000 731.000000 468.150000 ;
        RECT 721.000000 471.850000 731.000000 472.150000 ;
        RECT 710.000000 455.850000 715.000000 456.150000 ;
        RECT 710.000000 459.850000 715.000000 460.150000 ;
        RECT 710.000000 463.850000 715.000000 464.150000 ;
        RECT 710.000000 467.850000 715.000000 468.150000 ;
        RECT 710.000000 471.850000 715.000000 472.150000 ;
        RECT 721.000000 487.850000 731.000000 488.150000 ;
        RECT 721.000000 483.850000 731.000000 484.150000 ;
        RECT 721.000000 479.850000 731.000000 480.150000 ;
        RECT 721.000000 475.850000 731.000000 476.150000 ;
        RECT 710.000000 487.850000 715.000000 488.150000 ;
        RECT 710.000000 483.850000 715.000000 484.150000 ;
        RECT 710.000000 475.850000 715.000000 476.150000 ;
        RECT 710.000000 479.850000 715.000000 480.150000 ;
        RECT 810.000000 379.850000 815.000000 380.150000 ;
        RECT 760.000000 379.850000 765.000000 380.150000 ;
        RECT 760.000000 343.850000 765.000000 344.150000 ;
        RECT 760.000000 347.850000 765.000000 348.150000 ;
        RECT 760.000000 351.850000 765.000000 352.150000 ;
        RECT 760.000000 355.850000 765.000000 356.150000 ;
        RECT 760.000000 359.850000 765.000000 360.150000 ;
        RECT 760.000000 375.850000 765.000000 376.150000 ;
        RECT 760.000000 371.850000 765.000000 372.150000 ;
        RECT 760.000000 367.850000 765.000000 368.150000 ;
        RECT 760.000000 363.850000 765.000000 364.150000 ;
        RECT 810.000000 343.850000 815.000000 344.150000 ;
        RECT 810.000000 347.850000 815.000000 348.150000 ;
        RECT 810.000000 351.850000 815.000000 352.150000 ;
        RECT 810.000000 359.850000 815.000000 360.150000 ;
        RECT 810.000000 355.850000 815.000000 356.150000 ;
        RECT 810.000000 363.850000 815.000000 364.150000 ;
        RECT 810.000000 367.850000 815.000000 368.150000 ;
        RECT 810.000000 375.850000 815.000000 376.150000 ;
        RECT 810.000000 371.850000 815.000000 372.150000 ;
        RECT 760.000000 383.850000 765.000000 384.150000 ;
        RECT 760.000000 387.850000 765.000000 388.150000 ;
        RECT 760.000000 391.850000 765.000000 392.150000 ;
        RECT 760.000000 395.850000 765.000000 396.150000 ;
        RECT 760.000000 407.850000 765.000000 408.150000 ;
        RECT 760.000000 399.850000 765.000000 400.150000 ;
        RECT 760.000000 403.850000 765.000000 404.150000 ;
        RECT 760.000000 411.850000 765.000000 412.150000 ;
        RECT 760.000000 415.850000 765.000000 416.150000 ;
        RECT 810.000000 387.850000 815.000000 388.150000 ;
        RECT 810.000000 383.850000 815.000000 384.150000 ;
        RECT 810.000000 391.850000 815.000000 392.150000 ;
        RECT 810.000000 395.850000 815.000000 396.150000 ;
        RECT 810.000000 407.850000 815.000000 408.150000 ;
        RECT 810.000000 399.850000 815.000000 400.150000 ;
        RECT 810.000000 403.850000 815.000000 404.150000 ;
        RECT 810.000000 415.850000 815.000000 416.150000 ;
        RECT 810.000000 411.850000 815.000000 412.150000 ;
        RECT 860.000000 379.850000 865.000000 380.150000 ;
        RECT 860.000000 359.850000 865.000000 360.150000 ;
        RECT 860.000000 355.850000 865.000000 356.150000 ;
        RECT 860.000000 351.850000 865.000000 352.150000 ;
        RECT 860.000000 347.850000 865.000000 348.150000 ;
        RECT 860.000000 343.850000 865.000000 344.150000 ;
        RECT 860.000000 375.850000 865.000000 376.150000 ;
        RECT 860.000000 371.850000 865.000000 372.150000 ;
        RECT 860.000000 367.850000 865.000000 368.150000 ;
        RECT 860.000000 363.850000 865.000000 364.150000 ;
        RECT 860.000000 383.850000 865.000000 384.150000 ;
        RECT 860.000000 387.850000 865.000000 388.150000 ;
        RECT 860.000000 391.850000 865.000000 392.150000 ;
        RECT 860.000000 395.850000 865.000000 396.150000 ;
        RECT 860.000000 407.850000 865.000000 408.150000 ;
        RECT 860.000000 403.850000 865.000000 404.150000 ;
        RECT 860.000000 399.850000 865.000000 400.150000 ;
        RECT 860.000000 415.850000 865.000000 416.150000 ;
        RECT 860.000000 411.850000 865.000000 412.150000 ;
        RECT 760.000000 419.850000 765.000000 420.150000 ;
        RECT 760.000000 423.850000 765.000000 424.150000 ;
        RECT 760.000000 427.850000 765.000000 428.150000 ;
        RECT 760.000000 431.850000 765.000000 432.150000 ;
        RECT 760.000000 435.850000 765.000000 436.150000 ;
        RECT 760.000000 439.850000 765.000000 440.150000 ;
        RECT 760.000000 443.850000 765.000000 444.150000 ;
        RECT 810.000000 419.850000 815.000000 420.150000 ;
        RECT 810.000000 423.850000 815.000000 424.150000 ;
        RECT 810.000000 427.850000 815.000000 428.150000 ;
        RECT 810.000000 431.850000 815.000000 432.150000 ;
        RECT 810.000000 435.850000 815.000000 436.150000 ;
        RECT 810.000000 439.850000 815.000000 440.150000 ;
        RECT 810.000000 443.850000 815.000000 444.150000 ;
        RECT 860.000000 419.850000 865.000000 420.150000 ;
        RECT 860.000000 423.850000 865.000000 424.150000 ;
        RECT 860.000000 427.850000 865.000000 428.150000 ;
        RECT 860.000000 431.850000 865.000000 432.150000 ;
        RECT 860.000000 443.850000 865.000000 444.150000 ;
        RECT 860.000000 439.850000 865.000000 440.150000 ;
        RECT 860.000000 435.850000 865.000000 436.150000 ;
        RECT 610.000000 503.850000 615.000000 504.150000 ;
        RECT 610.000000 499.850000 615.000000 500.150000 ;
        RECT 610.000000 491.850000 615.000000 492.150000 ;
        RECT 610.000000 495.850000 615.000000 496.150000 ;
        RECT 660.000000 495.850000 665.000000 496.150000 ;
        RECT 660.000000 491.850000 665.000000 492.150000 ;
        RECT 660.000000 499.850000 665.000000 500.150000 ;
        RECT 660.000000 503.850000 665.000000 504.150000 ;
        RECT 710.000000 503.850000 715.000000 504.150000 ;
        RECT 710.000000 499.850000 715.000000 500.150000 ;
        RECT 710.000000 495.850000 715.000000 496.150000 ;
        RECT 710.000000 491.850000 715.000000 492.150000 ;
        RECT 960.000000 379.850000 965.000000 380.150000 ;
        RECT 960.000000 343.850000 965.000000 344.150000 ;
        RECT 960.000000 347.850000 965.000000 348.150000 ;
        RECT 960.000000 351.850000 965.000000 352.150000 ;
        RECT 960.000000 355.850000 965.000000 356.150000 ;
        RECT 960.000000 359.850000 965.000000 360.150000 ;
        RECT 960.000000 375.850000 965.000000 376.150000 ;
        RECT 960.000000 371.850000 965.000000 372.150000 ;
        RECT 960.000000 367.850000 965.000000 368.150000 ;
        RECT 960.000000 363.850000 965.000000 364.150000 ;
        RECT 960.000000 383.850000 965.000000 384.150000 ;
        RECT 960.000000 387.850000 965.000000 388.150000 ;
        RECT 960.000000 391.850000 965.000000 392.150000 ;
        RECT 960.000000 395.850000 965.000000 396.150000 ;
        RECT 960.000000 407.850000 965.000000 408.150000 ;
        RECT 960.000000 399.850000 965.000000 400.150000 ;
        RECT 960.000000 403.850000 965.000000 404.150000 ;
        RECT 960.000000 411.850000 965.000000 412.150000 ;
        RECT 960.000000 415.850000 965.000000 416.150000 ;
        RECT 910.000000 379.850000 915.000000 380.150000 ;
        RECT 910.000000 343.850000 915.000000 344.150000 ;
        RECT 910.000000 347.850000 915.000000 348.150000 ;
        RECT 910.000000 351.850000 915.000000 352.150000 ;
        RECT 910.000000 355.850000 915.000000 356.150000 ;
        RECT 910.000000 359.850000 915.000000 360.150000 ;
        RECT 910.000000 375.850000 915.000000 376.150000 ;
        RECT 910.000000 371.850000 915.000000 372.150000 ;
        RECT 910.000000 367.850000 915.000000 368.150000 ;
        RECT 910.000000 363.850000 915.000000 364.150000 ;
        RECT 910.000000 383.850000 915.000000 384.150000 ;
        RECT 910.000000 387.850000 915.000000 388.150000 ;
        RECT 910.000000 391.850000 915.000000 392.150000 ;
        RECT 910.000000 395.850000 915.000000 396.150000 ;
        RECT 910.000000 407.850000 915.000000 408.150000 ;
        RECT 910.000000 399.850000 915.000000 400.150000 ;
        RECT 910.000000 403.850000 915.000000 404.150000 ;
        RECT 910.000000 411.850000 915.000000 412.150000 ;
        RECT 910.000000 415.850000 915.000000 416.150000 ;
        RECT 1010.000000 379.850000 1015.000000 380.150000 ;
        RECT 1010.000000 343.850000 1015.000000 344.150000 ;
        RECT 1010.000000 347.850000 1015.000000 348.150000 ;
        RECT 1010.000000 351.850000 1015.000000 352.150000 ;
        RECT 1010.000000 359.850000 1015.000000 360.150000 ;
        RECT 1010.000000 355.850000 1015.000000 356.150000 ;
        RECT 1010.000000 363.850000 1015.000000 364.150000 ;
        RECT 1010.000000 367.850000 1015.000000 368.150000 ;
        RECT 1010.000000 375.850000 1015.000000 376.150000 ;
        RECT 1010.000000 371.850000 1015.000000 372.150000 ;
        RECT 1010.000000 387.850000 1015.000000 388.150000 ;
        RECT 1010.000000 383.850000 1015.000000 384.150000 ;
        RECT 1010.000000 391.850000 1015.000000 392.150000 ;
        RECT 1010.000000 395.850000 1015.000000 396.150000 ;
        RECT 1010.000000 407.850000 1015.000000 408.150000 ;
        RECT 1010.000000 403.850000 1015.000000 404.150000 ;
        RECT 1010.000000 399.850000 1015.000000 400.150000 ;
        RECT 1010.000000 415.850000 1015.000000 416.150000 ;
        RECT 1010.000000 411.850000 1015.000000 412.150000 ;
        RECT 960.000000 431.850000 965.000000 432.150000 ;
        RECT 960.000000 427.850000 965.000000 428.150000 ;
        RECT 960.000000 423.850000 965.000000 424.150000 ;
        RECT 960.000000 419.850000 965.000000 420.150000 ;
        RECT 960.000000 443.850000 965.000000 444.150000 ;
        RECT 960.000000 439.850000 965.000000 440.150000 ;
        RECT 960.000000 435.850000 965.000000 436.150000 ;
        RECT 910.000000 419.850000 915.000000 420.150000 ;
        RECT 910.000000 423.850000 915.000000 424.150000 ;
        RECT 910.000000 427.850000 915.000000 428.150000 ;
        RECT 910.000000 431.850000 915.000000 432.150000 ;
        RECT 910.000000 435.850000 915.000000 436.150000 ;
        RECT 910.000000 439.850000 915.000000 440.150000 ;
        RECT 910.000000 443.850000 915.000000 444.150000 ;
        RECT 1010.000000 419.850000 1015.000000 420.150000 ;
        RECT 1010.000000 423.850000 1015.000000 424.150000 ;
        RECT 1010.000000 427.850000 1015.000000 428.150000 ;
        RECT 1010.000000 431.850000 1015.000000 432.150000 ;
        RECT 1010.000000 439.850000 1015.000000 440.150000 ;
        RECT 1010.000000 435.850000 1015.000000 436.150000 ;
        RECT 1010.000000 443.850000 1015.000000 444.150000 ;
        RECT 1110.000000 379.850000 1115.000000 380.150000 ;
        RECT 1110.000000 343.850000 1115.000000 344.150000 ;
        RECT 1110.000000 347.850000 1115.000000 348.150000 ;
        RECT 1110.000000 351.850000 1115.000000 352.150000 ;
        RECT 1110.000000 355.850000 1115.000000 356.150000 ;
        RECT 1110.000000 359.850000 1115.000000 360.150000 ;
        RECT 1110.000000 375.850000 1115.000000 376.150000 ;
        RECT 1110.000000 371.850000 1115.000000 372.150000 ;
        RECT 1110.000000 367.850000 1115.000000 368.150000 ;
        RECT 1110.000000 363.850000 1115.000000 364.150000 ;
        RECT 1110.000000 383.850000 1115.000000 384.150000 ;
        RECT 1110.000000 387.850000 1115.000000 388.150000 ;
        RECT 1110.000000 391.850000 1115.000000 392.150000 ;
        RECT 1110.000000 395.850000 1115.000000 396.150000 ;
        RECT 1110.000000 407.850000 1115.000000 408.150000 ;
        RECT 1110.000000 399.850000 1115.000000 400.150000 ;
        RECT 1110.000000 403.850000 1115.000000 404.150000 ;
        RECT 1110.000000 411.850000 1115.000000 412.150000 ;
        RECT 1110.000000 415.850000 1115.000000 416.150000 ;
        RECT 1060.000000 379.850000 1065.000000 380.150000 ;
        RECT 1060.000000 343.850000 1065.000000 344.150000 ;
        RECT 1060.000000 347.850000 1065.000000 348.150000 ;
        RECT 1060.000000 351.850000 1065.000000 352.150000 ;
        RECT 1060.000000 355.850000 1065.000000 356.150000 ;
        RECT 1060.000000 359.850000 1065.000000 360.150000 ;
        RECT 1060.000000 375.850000 1065.000000 376.150000 ;
        RECT 1060.000000 371.850000 1065.000000 372.150000 ;
        RECT 1060.000000 367.850000 1065.000000 368.150000 ;
        RECT 1060.000000 363.850000 1065.000000 364.150000 ;
        RECT 1060.000000 395.850000 1065.000000 396.150000 ;
        RECT 1060.000000 391.850000 1065.000000 392.150000 ;
        RECT 1060.000000 387.850000 1065.000000 388.150000 ;
        RECT 1060.000000 383.850000 1065.000000 384.150000 ;
        RECT 1060.000000 407.850000 1065.000000 408.150000 ;
        RECT 1060.000000 403.850000 1065.000000 404.150000 ;
        RECT 1060.000000 399.850000 1065.000000 400.150000 ;
        RECT 1060.000000 411.850000 1065.000000 412.150000 ;
        RECT 1060.000000 415.850000 1065.000000 416.150000 ;
        RECT 1158.000000 379.850000 1168.000000 380.150000 ;
        RECT 1158.000000 343.850000 1168.000000 344.150000 ;
        RECT 1158.000000 347.850000 1168.000000 348.150000 ;
        RECT 1158.000000 351.850000 1168.000000 352.150000 ;
        RECT 1158.000000 355.850000 1168.000000 356.150000 ;
        RECT 1158.000000 359.850000 1168.000000 360.150000 ;
        RECT 1158.000000 375.850000 1168.000000 376.150000 ;
        RECT 1158.000000 371.850000 1168.000000 372.150000 ;
        RECT 1158.000000 367.850000 1168.000000 368.150000 ;
        RECT 1158.000000 363.850000 1168.000000 364.150000 ;
        RECT 1158.000000 395.850000 1168.000000 396.150000 ;
        RECT 1158.000000 391.850000 1168.000000 392.150000 ;
        RECT 1158.000000 387.850000 1168.000000 388.150000 ;
        RECT 1158.000000 383.850000 1168.000000 384.150000 ;
        RECT 1158.000000 407.850000 1168.000000 408.150000 ;
        RECT 1158.000000 399.850000 1168.000000 400.150000 ;
        RECT 1158.000000 403.850000 1168.000000 404.150000 ;
        RECT 1158.000000 411.850000 1168.000000 412.150000 ;
        RECT 1158.000000 415.850000 1168.000000 416.150000 ;
        RECT 1110.000000 431.850000 1115.000000 432.150000 ;
        RECT 1110.000000 427.850000 1115.000000 428.150000 ;
        RECT 1110.000000 423.850000 1115.000000 424.150000 ;
        RECT 1110.000000 419.850000 1115.000000 420.150000 ;
        RECT 1110.000000 443.850000 1115.000000 444.150000 ;
        RECT 1110.000000 439.850000 1115.000000 440.150000 ;
        RECT 1110.000000 435.850000 1115.000000 436.150000 ;
        RECT 1060.000000 419.850000 1065.000000 420.150000 ;
        RECT 1060.000000 423.850000 1065.000000 424.150000 ;
        RECT 1060.000000 431.850000 1065.000000 432.150000 ;
        RECT 1060.000000 427.850000 1065.000000 428.150000 ;
        RECT 1060.000000 435.850000 1065.000000 436.150000 ;
        RECT 1060.000000 439.850000 1065.000000 440.150000 ;
        RECT 1060.000000 443.850000 1065.000000 444.150000 ;
        RECT 1158.000000 427.850000 1168.000000 428.150000 ;
        RECT 1158.000000 423.850000 1168.000000 424.150000 ;
        RECT 1158.000000 419.850000 1168.000000 420.150000 ;
        RECT 1160.000000 431.850000 1165.000000 432.150000 ;
        RECT 1160.000000 435.850000 1165.000000 436.150000 ;
        RECT 1160.000000 439.850000 1165.000000 440.150000 ;
        RECT 1160.000000 443.850000 1165.000000 444.150000 ;
        RECT 1160.000000 447.850000 1165.000000 448.150000 ;
        RECT 1160.000000 451.850000 1165.000000 452.150000 ;
        RECT 1160.000000 459.850000 1165.000000 460.150000 ;
        RECT 1160.000000 455.850000 1165.000000 456.150000 ;
        RECT 1160.000000 463.850000 1165.000000 464.150000 ;
        RECT 1160.000000 467.850000 1165.000000 468.150000 ;
        RECT 1160.000000 471.850000 1165.000000 472.150000 ;
        RECT 1160.000000 479.850000 1165.000000 480.150000 ;
        RECT 1160.000000 475.850000 1165.000000 476.150000 ;
        RECT 1160.000000 487.850000 1165.000000 488.150000 ;
        RECT 1160.000000 483.850000 1165.000000 484.150000 ;
        RECT 1160.000000 491.850000 1165.000000 492.150000 ;
        RECT 1160.000000 495.850000 1165.000000 496.150000 ;
        RECT 1160.000000 499.850000 1165.000000 500.150000 ;
        RECT 1160.000000 507.850000 1165.000000 508.150000 ;
        RECT 1160.000000 503.850000 1165.000000 504.150000 ;
        RECT 1160.000000 511.850000 1165.000000 512.150000 ;
        RECT 1160.000000 515.850000 1165.000000 516.150000 ;
        RECT 1160.000000 519.850000 1165.000000 520.150000 ;
        RECT 1160.000000 523.850000 1165.000000 524.150000 ;
        RECT 1160.000000 527.850000 1165.000000 528.150000 ;
        RECT 1160.000000 535.850000 1165.000000 536.150000 ;
        RECT 1160.000000 531.850000 1165.000000 532.150000 ;
        RECT 1160.000000 539.850000 1165.000000 540.150000 ;
        RECT 1160.000000 543.850000 1165.000000 544.150000 ;
        RECT 1160.000000 555.850000 1165.000000 556.150000 ;
        RECT 1160.000000 551.850000 1165.000000 552.150000 ;
        RECT 1160.000000 547.850000 1165.000000 548.150000 ;
        RECT 1160.000000 563.850000 1165.000000 564.150000 ;
        RECT 1160.000000 559.850000 1165.000000 560.150000 ;
        RECT 1160.000000 583.850000 1165.000000 584.150000 ;
        RECT 1160.000000 567.850000 1165.000000 568.150000 ;
        RECT 1160.000000 571.850000 1165.000000 572.150000 ;
        RECT 1160.000000 579.850000 1165.000000 580.150000 ;
        RECT 1160.000000 575.850000 1165.000000 576.150000 ;
        RECT 1160.000000 591.850000 1165.000000 592.150000 ;
        RECT 1160.000000 587.850000 1165.000000 588.150000 ;
        RECT 1160.000000 595.850000 1165.000000 596.150000 ;
        RECT 1160.000000 599.850000 1165.000000 600.150000 ;
        RECT 1160.000000 607.850000 1165.000000 608.150000 ;
        RECT 1160.000000 603.850000 1165.000000 604.150000 ;
        RECT 1160.000000 611.850000 1165.000000 612.150000 ;
        RECT 1160.000000 615.850000 1165.000000 616.150000 ;
        RECT 1160.000000 619.850000 1165.000000 620.150000 ;
        RECT 1160.000000 623.850000 1165.000000 624.150000 ;
        RECT 1160.000000 627.850000 1165.000000 628.150000 ;
        RECT 1160.000000 635.850000 1165.000000 636.150000 ;
        RECT 1160.000000 631.850000 1165.000000 632.150000 ;
        RECT 610.000000 659.850000 615.000000 660.150000 ;
        RECT 610.000000 663.850000 615.000000 664.150000 ;
        RECT 610.000000 667.850000 615.000000 668.150000 ;
        RECT 610.000000 671.850000 615.000000 672.150000 ;
        RECT 610.000000 675.850000 615.000000 676.150000 ;
        RECT 660.000000 663.850000 665.000000 664.150000 ;
        RECT 660.000000 659.850000 665.000000 660.150000 ;
        RECT 660.000000 667.850000 665.000000 668.150000 ;
        RECT 660.000000 671.850000 665.000000 672.150000 ;
        RECT 660.000000 675.850000 665.000000 676.150000 ;
        RECT 610.000000 683.850000 615.000000 684.150000 ;
        RECT 610.000000 679.850000 615.000000 680.150000 ;
        RECT 660.000000 683.850000 665.000000 684.150000 ;
        RECT 660.000000 679.850000 665.000000 680.150000 ;
        RECT 1160.000000 639.850000 1165.000000 640.150000 ;
        RECT 1160.000000 643.850000 1165.000000 644.150000 ;
        RECT 1160.000000 647.850000 1165.000000 648.150000 ;
        RECT 1160.000000 655.850000 1165.000000 656.150000 ;
        RECT 1160.000000 651.850000 1165.000000 652.150000 ;
        RECT 1160.000000 663.850000 1165.000000 664.150000 ;
        RECT 1160.000000 659.850000 1165.000000 660.150000 ;
        RECT 1160.000000 667.850000 1165.000000 668.150000 ;
        RECT 1160.000000 671.850000 1165.000000 672.150000 ;
        RECT 1160.000000 675.850000 1165.000000 676.150000 ;
        RECT 1160.000000 683.850000 1165.000000 684.150000 ;
        RECT 1160.000000 679.850000 1165.000000 680.150000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  OBS
    LAYER OVERLAP ;
      RECT 0.000000 656.000000 670.000000 686.000000 ;
      RECT 0.000000 506.000000 399.000000 656.000000 ;
      RECT 1139.000000 446.000000 1186.000000 686.000000 ;
      RECT 0.000000 446.000000 749.000000 506.000000 ;
      RECT 0.000000 0.000000 1186.000000 446.000000 ;
    LAYER M1 ;
      RECT 0.000000 656.000000 670.000000 686.000000 ;
      RECT 0.000000 506.000000 399.000000 656.000000 ;
      RECT 1139.000000 446.000000 1186.000000 686.000000 ;
      RECT 0.000000 446.000000 749.000000 506.000000 ;
      RECT 0.000000 0.000000 1186.000000 446.000000 ;
    LAYER M2 ;
      RECT 1139.000000 685.650000 1186.000000 686.000000 ;
      RECT 647.765000 685.650000 670.000000 686.000000 ;
      RECT 561.965000 685.650000 624.430000 686.000000 ;
      RECT 556.285000 685.650000 558.865000 686.000000 ;
      RECT 476.165000 685.650000 538.630000 686.000000 ;
      RECT 455.930000 685.650000 463.425000 686.000000 ;
      RECT 390.365000 685.650000 452.830000 686.000000 ;
      RECT 304.565000 685.650000 367.030000 686.000000 ;
      RECT 647.765000 683.980000 658.500000 685.650000 ;
      RECT 642.085000 683.980000 644.665000 686.000000 ;
      RECT 638.125000 683.980000 638.985000 686.000000 ;
      RECT 627.530000 683.980000 635.025000 686.000000 ;
      RECT 616.500000 683.980000 624.430000 685.650000 ;
      RECT 556.285000 683.980000 558.500000 685.650000 ;
      RECT 552.325000 683.980000 553.185000 686.000000 ;
      RECT 541.730000 683.980000 549.225000 686.000000 ;
      RECT 516.500000 683.980000 538.630000 685.650000 ;
      RECT 476.165000 683.980000 508.500000 685.650000 ;
      RECT 470.485000 683.980000 473.065000 686.000000 ;
      RECT 466.525000 683.980000 467.385000 686.000000 ;
      RECT 455.930000 683.980000 458.500000 685.650000 ;
      RECT 416.500000 683.980000 452.830000 685.650000 ;
      RECT 390.365000 683.980000 408.500000 685.650000 ;
      RECT 384.685000 683.980000 387.265000 686.000000 ;
      RECT 380.725000 683.980000 381.585000 686.000000 ;
      RECT 370.130000 683.980000 377.625000 686.000000 ;
      RECT 366.500000 683.980000 367.030000 685.650000 ;
      RECT 304.565000 683.980000 308.500000 685.650000 ;
      RECT 298.885000 683.980000 301.465000 686.000000 ;
      RECT 294.925000 683.980000 295.785000 686.000000 ;
      RECT 284.330000 683.980000 291.825000 686.000000 ;
      RECT 218.765000 683.980000 281.230000 686.000000 ;
      RECT 213.085000 683.980000 215.665000 686.000000 ;
      RECT 209.125000 683.980000 209.985000 686.000000 ;
      RECT 198.530000 683.980000 206.025000 686.000000 ;
      RECT 132.965000 683.980000 195.430000 686.000000 ;
      RECT 127.285000 683.980000 129.865000 686.000000 ;
      RECT 123.325000 683.980000 124.185000 686.000000 ;
      RECT 112.730000 683.980000 120.225000 686.000000 ;
      RECT 47.165000 683.980000 109.630000 686.000000 ;
      RECT 41.485000 683.980000 44.065000 686.000000 ;
      RECT 37.525000 683.980000 38.385000 686.000000 ;
      RECT 26.930000 683.980000 34.425000 686.000000 ;
      RECT 0.000000 683.980000 23.830000 686.000000 ;
      RECT 1139.000000 683.650000 1158.500000 685.650000 ;
      RECT 616.500000 683.650000 658.500000 683.980000 ;
      RECT 566.500000 683.650000 608.500000 685.650000 ;
      RECT 516.500000 683.650000 558.500000 683.980000 ;
      RECT 466.500000 683.650000 508.500000 683.980000 ;
      RECT 416.500000 683.650000 458.500000 683.980000 ;
      RECT 366.500000 683.650000 408.500000 683.980000 ;
      RECT 316.500000 683.650000 358.500000 685.650000 ;
      RECT 0.000000 683.650000 308.500000 683.980000 ;
      RECT 1166.500000 682.350000 1186.000000 685.650000 ;
      RECT 1157.500000 682.350000 1158.500000 683.650000 ;
      RECT 666.500000 682.350000 670.000000 685.650000 ;
      RECT 657.500000 682.350000 658.500000 683.650000 ;
      RECT 616.500000 682.350000 649.500000 683.650000 ;
      RECT 607.500000 682.350000 608.500000 683.650000 ;
      RECT 566.500000 682.350000 599.500000 683.650000 ;
      RECT 557.500000 682.350000 558.500000 683.650000 ;
      RECT 516.500000 682.350000 549.500000 683.650000 ;
      RECT 507.500000 682.350000 508.500000 683.650000 ;
      RECT 466.500000 682.350000 499.500000 683.650000 ;
      RECT 457.500000 682.350000 458.500000 683.650000 ;
      RECT 416.500000 682.350000 449.500000 683.650000 ;
      RECT 407.500000 682.350000 408.500000 683.650000 ;
      RECT 366.500000 682.350000 383.500000 683.650000 ;
      RECT 357.500000 682.350000 358.500000 683.650000 ;
      RECT 316.500000 682.350000 349.500000 683.650000 ;
      RECT 307.500000 682.350000 308.500000 683.650000 ;
      RECT 1157.500000 681.650000 1186.000000 682.350000 ;
      RECT 657.500000 681.650000 670.000000 682.350000 ;
      RECT 607.500000 681.650000 649.500000 682.350000 ;
      RECT 557.500000 681.650000 599.500000 682.350000 ;
      RECT 507.500000 681.650000 549.500000 682.350000 ;
      RECT 457.500000 681.650000 499.500000 682.350000 ;
      RECT 407.500000 681.650000 449.500000 682.350000 ;
      RECT 357.500000 681.650000 383.500000 682.350000 ;
      RECT 307.500000 681.650000 349.500000 682.350000 ;
      RECT 1157.500000 680.350000 1158.500000 681.650000 ;
      RECT 1139.000000 680.350000 1149.500000 683.650000 ;
      RECT 657.500000 680.350000 658.500000 681.650000 ;
      RECT 616.500000 680.350000 649.500000 681.650000 ;
      RECT 607.500000 680.350000 608.500000 681.650000 ;
      RECT 566.500000 680.350000 599.500000 681.650000 ;
      RECT 557.500000 680.350000 558.500000 681.650000 ;
      RECT 516.500000 680.350000 549.500000 681.650000 ;
      RECT 507.500000 680.350000 508.500000 681.650000 ;
      RECT 466.500000 680.350000 499.500000 681.650000 ;
      RECT 457.500000 680.350000 458.500000 681.650000 ;
      RECT 416.500000 680.350000 449.500000 681.650000 ;
      RECT 407.500000 680.350000 408.500000 681.650000 ;
      RECT 396.500000 680.350000 399.500000 683.650000 ;
      RECT 366.500000 680.350000 383.500000 681.650000 ;
      RECT 357.500000 680.350000 358.500000 681.650000 ;
      RECT 316.500000 680.350000 349.500000 681.650000 ;
      RECT 307.500000 680.350000 308.500000 681.650000 ;
      RECT 0.000000 680.350000 299.500000 683.650000 ;
      RECT 1139.000000 679.650000 1158.500000 680.350000 ;
      RECT 616.500000 679.650000 658.500000 680.350000 ;
      RECT 566.500000 679.650000 608.500000 680.350000 ;
      RECT 516.500000 679.650000 558.500000 680.350000 ;
      RECT 466.500000 679.650000 508.500000 680.350000 ;
      RECT 416.500000 679.650000 458.500000 680.350000 ;
      RECT 366.500000 679.650000 408.500000 680.350000 ;
      RECT 316.500000 679.650000 358.500000 680.350000 ;
      RECT 0.000000 679.650000 308.500000 680.350000 ;
      RECT 1166.500000 678.350000 1186.000000 681.650000 ;
      RECT 1157.500000 678.350000 1158.500000 679.650000 ;
      RECT 666.500000 678.350000 670.000000 681.650000 ;
      RECT 657.500000 678.350000 658.500000 679.650000 ;
      RECT 616.500000 678.350000 649.500000 679.650000 ;
      RECT 607.500000 678.350000 608.500000 679.650000 ;
      RECT 566.500000 678.350000 599.500000 679.650000 ;
      RECT 557.500000 678.350000 558.500000 679.650000 ;
      RECT 516.500000 678.350000 549.500000 679.650000 ;
      RECT 507.500000 678.350000 508.500000 679.650000 ;
      RECT 466.500000 678.350000 499.500000 679.650000 ;
      RECT 457.500000 678.350000 458.500000 679.650000 ;
      RECT 416.500000 678.350000 449.500000 679.650000 ;
      RECT 407.500000 678.350000 408.500000 679.650000 ;
      RECT 366.500000 678.350000 383.500000 679.650000 ;
      RECT 357.500000 678.350000 358.500000 679.650000 ;
      RECT 316.500000 678.350000 349.500000 679.650000 ;
      RECT 307.500000 678.350000 308.500000 679.650000 ;
      RECT 1157.500000 677.650000 1186.000000 678.350000 ;
      RECT 657.500000 677.650000 670.000000 678.350000 ;
      RECT 607.500000 677.650000 649.500000 678.350000 ;
      RECT 557.500000 677.650000 599.500000 678.350000 ;
      RECT 507.500000 677.650000 549.500000 678.350000 ;
      RECT 457.500000 677.650000 499.500000 678.350000 ;
      RECT 407.500000 677.650000 449.500000 678.350000 ;
      RECT 357.500000 677.650000 383.500000 678.350000 ;
      RECT 1157.500000 676.350000 1158.500000 677.650000 ;
      RECT 1139.000000 676.350000 1149.500000 679.650000 ;
      RECT 657.500000 676.350000 658.500000 677.650000 ;
      RECT 616.500000 676.350000 649.500000 677.650000 ;
      RECT 607.500000 676.350000 608.500000 677.650000 ;
      RECT 566.500000 676.350000 599.500000 677.650000 ;
      RECT 557.500000 676.350000 558.500000 677.650000 ;
      RECT 516.500000 676.350000 549.500000 677.650000 ;
      RECT 507.500000 676.350000 508.500000 677.650000 ;
      RECT 466.500000 676.350000 499.500000 677.650000 ;
      RECT 457.500000 676.350000 458.500000 677.650000 ;
      RECT 416.500000 676.350000 449.500000 677.650000 ;
      RECT 407.500000 676.350000 408.500000 677.650000 ;
      RECT 396.500000 676.350000 399.500000 679.650000 ;
      RECT 366.500000 676.350000 383.500000 677.650000 ;
      RECT 357.500000 676.350000 358.500000 677.650000 ;
      RECT 307.500000 676.350000 349.500000 678.350000 ;
      RECT 0.000000 676.350000 299.500000 679.650000 ;
      RECT 1139.000000 675.650000 1158.500000 676.350000 ;
      RECT 616.500000 675.650000 658.500000 676.350000 ;
      RECT 566.500000 675.650000 608.500000 676.350000 ;
      RECT 516.500000 675.650000 558.500000 676.350000 ;
      RECT 466.500000 675.650000 508.500000 676.350000 ;
      RECT 416.500000 675.650000 458.500000 676.350000 ;
      RECT 366.500000 675.650000 408.500000 676.350000 ;
      RECT 0.000000 675.650000 358.500000 676.350000 ;
      RECT 1166.500000 674.350000 1186.000000 677.650000 ;
      RECT 1157.500000 674.350000 1158.500000 675.650000 ;
      RECT 666.500000 674.350000 670.000000 677.650000 ;
      RECT 657.500000 674.350000 658.500000 675.650000 ;
      RECT 616.500000 674.350000 649.500000 675.650000 ;
      RECT 607.500000 674.350000 608.500000 675.650000 ;
      RECT 566.500000 674.350000 599.500000 675.650000 ;
      RECT 557.500000 674.350000 558.500000 675.650000 ;
      RECT 516.500000 674.350000 549.500000 675.650000 ;
      RECT 507.500000 674.350000 508.500000 675.650000 ;
      RECT 466.500000 674.350000 499.500000 675.650000 ;
      RECT 457.500000 674.350000 458.500000 675.650000 ;
      RECT 416.500000 674.350000 449.500000 675.650000 ;
      RECT 407.500000 674.350000 408.500000 675.650000 ;
      RECT 366.500000 674.350000 383.500000 675.650000 ;
      RECT 357.500000 674.350000 358.500000 675.650000 ;
      RECT 1157.500000 673.650000 1186.000000 674.350000 ;
      RECT 657.500000 673.650000 670.000000 674.350000 ;
      RECT 607.500000 673.650000 649.500000 674.350000 ;
      RECT 557.500000 673.650000 599.500000 674.350000 ;
      RECT 507.500000 673.650000 549.500000 674.350000 ;
      RECT 457.500000 673.650000 499.500000 674.350000 ;
      RECT 407.500000 673.650000 449.500000 674.350000 ;
      RECT 357.500000 673.650000 383.500000 674.350000 ;
      RECT 1157.500000 672.350000 1158.500000 673.650000 ;
      RECT 1139.000000 672.350000 1149.500000 675.650000 ;
      RECT 657.500000 672.350000 658.500000 673.650000 ;
      RECT 616.500000 672.350000 649.500000 673.650000 ;
      RECT 607.500000 672.350000 608.500000 673.650000 ;
      RECT 566.500000 672.350000 599.500000 673.650000 ;
      RECT 557.500000 672.350000 558.500000 673.650000 ;
      RECT 516.500000 672.350000 549.500000 673.650000 ;
      RECT 507.500000 672.350000 508.500000 673.650000 ;
      RECT 466.500000 672.350000 499.500000 673.650000 ;
      RECT 457.500000 672.350000 458.500000 673.650000 ;
      RECT 416.500000 672.350000 449.500000 673.650000 ;
      RECT 407.500000 672.350000 408.500000 673.650000 ;
      RECT 396.500000 672.350000 399.500000 675.650000 ;
      RECT 366.500000 672.350000 383.500000 673.650000 ;
      RECT 357.500000 672.350000 358.500000 673.650000 ;
      RECT 0.000000 672.350000 349.500000 675.650000 ;
      RECT 1139.000000 671.650000 1158.500000 672.350000 ;
      RECT 616.500000 671.650000 658.500000 672.350000 ;
      RECT 566.500000 671.650000 608.500000 672.350000 ;
      RECT 516.500000 671.650000 558.500000 672.350000 ;
      RECT 466.500000 671.650000 508.500000 672.350000 ;
      RECT 416.500000 671.650000 458.500000 672.350000 ;
      RECT 366.500000 671.650000 408.500000 672.350000 ;
      RECT 0.000000 671.650000 358.500000 672.350000 ;
      RECT 1166.500000 670.350000 1186.000000 673.650000 ;
      RECT 1157.500000 670.350000 1158.500000 671.650000 ;
      RECT 666.500000 670.350000 670.000000 673.650000 ;
      RECT 657.500000 670.350000 658.500000 671.650000 ;
      RECT 616.500000 670.350000 649.500000 671.650000 ;
      RECT 607.500000 670.350000 608.500000 671.650000 ;
      RECT 566.500000 670.350000 599.500000 671.650000 ;
      RECT 557.500000 670.350000 558.500000 671.650000 ;
      RECT 516.500000 670.350000 549.500000 671.650000 ;
      RECT 507.500000 670.350000 508.500000 671.650000 ;
      RECT 466.500000 670.350000 499.500000 671.650000 ;
      RECT 457.500000 670.350000 458.500000 671.650000 ;
      RECT 416.500000 670.350000 449.500000 671.650000 ;
      RECT 407.500000 670.350000 408.500000 671.650000 ;
      RECT 366.500000 670.350000 383.500000 671.650000 ;
      RECT 357.500000 670.350000 358.500000 671.650000 ;
      RECT 1157.500000 669.650000 1186.000000 670.350000 ;
      RECT 657.500000 669.650000 670.000000 670.350000 ;
      RECT 607.500000 669.650000 649.500000 670.350000 ;
      RECT 557.500000 669.650000 599.500000 670.350000 ;
      RECT 507.500000 669.650000 549.500000 670.350000 ;
      RECT 457.500000 669.650000 499.500000 670.350000 ;
      RECT 407.500000 669.650000 449.500000 670.350000 ;
      RECT 357.500000 669.650000 383.500000 670.350000 ;
      RECT 1157.500000 668.350000 1158.500000 669.650000 ;
      RECT 1139.000000 668.350000 1149.500000 671.650000 ;
      RECT 657.500000 668.350000 658.500000 669.650000 ;
      RECT 616.500000 668.350000 649.500000 669.650000 ;
      RECT 607.500000 668.350000 608.500000 669.650000 ;
      RECT 566.500000 668.350000 599.500000 669.650000 ;
      RECT 557.500000 668.350000 558.500000 669.650000 ;
      RECT 516.500000 668.350000 549.500000 669.650000 ;
      RECT 507.500000 668.350000 508.500000 669.650000 ;
      RECT 466.500000 668.350000 499.500000 669.650000 ;
      RECT 457.500000 668.350000 458.500000 669.650000 ;
      RECT 416.500000 668.350000 449.500000 669.650000 ;
      RECT 407.500000 668.350000 408.500000 669.650000 ;
      RECT 396.500000 668.350000 399.500000 671.650000 ;
      RECT 382.500000 668.350000 383.500000 669.650000 ;
      RECT 357.500000 668.350000 358.500000 669.650000 ;
      RECT 0.000000 668.350000 349.500000 671.650000 ;
      RECT 1139.000000 667.650000 1158.500000 668.350000 ;
      RECT 616.500000 667.650000 658.500000 668.350000 ;
      RECT 566.500000 667.650000 608.500000 668.350000 ;
      RECT 516.500000 667.650000 558.500000 668.350000 ;
      RECT 466.500000 667.650000 508.500000 668.350000 ;
      RECT 416.500000 667.650000 458.500000 668.350000 ;
      RECT 382.500000 667.650000 408.500000 668.350000 ;
      RECT 0.000000 667.650000 358.500000 668.350000 ;
      RECT 1166.500000 666.350000 1186.000000 669.650000 ;
      RECT 1157.500000 666.350000 1158.500000 667.650000 ;
      RECT 666.500000 666.350000 670.000000 669.650000 ;
      RECT 657.500000 666.350000 658.500000 667.650000 ;
      RECT 616.500000 666.350000 649.500000 667.650000 ;
      RECT 607.500000 666.350000 608.500000 667.650000 ;
      RECT 566.500000 666.350000 599.500000 667.650000 ;
      RECT 557.500000 666.350000 558.500000 667.650000 ;
      RECT 516.500000 666.350000 549.500000 667.650000 ;
      RECT 507.500000 666.350000 508.500000 667.650000 ;
      RECT 466.500000 666.350000 499.500000 667.650000 ;
      RECT 457.500000 666.350000 458.500000 667.650000 ;
      RECT 416.500000 666.350000 449.500000 667.650000 ;
      RECT 407.500000 666.350000 408.500000 667.650000 ;
      RECT 382.500000 666.350000 383.500000 667.650000 ;
      RECT 366.500000 666.350000 369.500000 669.650000 ;
      RECT 357.500000 666.350000 358.500000 667.650000 ;
      RECT 1157.500000 665.650000 1186.000000 666.350000 ;
      RECT 657.500000 665.650000 670.000000 666.350000 ;
      RECT 607.500000 665.650000 649.500000 666.350000 ;
      RECT 557.500000 665.650000 599.500000 666.350000 ;
      RECT 507.500000 665.650000 549.500000 666.350000 ;
      RECT 457.500000 665.650000 499.500000 666.350000 ;
      RECT 407.500000 665.650000 449.500000 666.350000 ;
      RECT 357.500000 665.650000 383.500000 666.350000 ;
      RECT 1157.500000 664.350000 1158.500000 665.650000 ;
      RECT 1139.000000 664.350000 1149.500000 667.650000 ;
      RECT 657.500000 664.350000 658.500000 665.650000 ;
      RECT 616.500000 664.350000 649.500000 665.650000 ;
      RECT 607.500000 664.350000 608.500000 665.650000 ;
      RECT 566.500000 664.350000 599.500000 665.650000 ;
      RECT 557.500000 664.350000 558.500000 665.650000 ;
      RECT 516.500000 664.350000 549.500000 665.650000 ;
      RECT 507.500000 664.350000 508.500000 665.650000 ;
      RECT 466.500000 664.350000 499.500000 665.650000 ;
      RECT 457.500000 664.350000 458.500000 665.650000 ;
      RECT 416.500000 664.350000 449.500000 665.650000 ;
      RECT 407.500000 664.350000 408.500000 665.650000 ;
      RECT 396.500000 664.350000 399.500000 667.650000 ;
      RECT 382.500000 664.350000 383.500000 665.650000 ;
      RECT 357.500000 664.350000 358.500000 665.650000 ;
      RECT 0.000000 664.350000 349.500000 667.650000 ;
      RECT 1139.000000 663.650000 1158.500000 664.350000 ;
      RECT 616.500000 663.650000 658.500000 664.350000 ;
      RECT 566.500000 663.650000 608.500000 664.350000 ;
      RECT 516.500000 663.650000 558.500000 664.350000 ;
      RECT 466.500000 663.650000 508.500000 664.350000 ;
      RECT 416.500000 663.650000 458.500000 664.350000 ;
      RECT 382.500000 663.650000 408.500000 664.350000 ;
      RECT 0.000000 663.650000 358.500000 664.350000 ;
      RECT 0.000000 663.170000 349.500000 663.650000 ;
      RECT 1166.500000 663.165000 1186.000000 665.650000 ;
      RECT 1166.500000 662.350000 1183.980000 663.165000 ;
      RECT 1157.500000 662.350000 1158.500000 663.650000 ;
      RECT 666.500000 662.350000 670.000000 665.650000 ;
      RECT 657.500000 662.350000 658.500000 663.650000 ;
      RECT 616.500000 662.350000 649.500000 663.650000 ;
      RECT 607.500000 662.350000 608.500000 663.650000 ;
      RECT 566.500000 662.350000 599.500000 663.650000 ;
      RECT 557.500000 662.350000 558.500000 663.650000 ;
      RECT 516.500000 662.350000 549.500000 663.650000 ;
      RECT 507.500000 662.350000 508.500000 663.650000 ;
      RECT 466.500000 662.350000 499.500000 663.650000 ;
      RECT 457.500000 662.350000 458.500000 663.650000 ;
      RECT 416.500000 662.350000 449.500000 663.650000 ;
      RECT 407.500000 662.350000 408.500000 663.650000 ;
      RECT 382.500000 662.350000 383.500000 663.650000 ;
      RECT 366.500000 662.350000 369.500000 665.650000 ;
      RECT 357.500000 662.350000 358.500000 663.650000 ;
      RECT 1157.500000 661.650000 1183.980000 662.350000 ;
      RECT 657.500000 661.650000 670.000000 662.350000 ;
      RECT 607.500000 661.650000 649.500000 662.350000 ;
      RECT 557.500000 661.650000 599.500000 662.350000 ;
      RECT 507.500000 661.650000 549.500000 662.350000 ;
      RECT 457.500000 661.650000 499.500000 662.350000 ;
      RECT 407.500000 661.650000 449.500000 662.350000 ;
      RECT 357.500000 661.650000 383.500000 662.350000 ;
      RECT 1157.500000 660.350000 1158.500000 661.650000 ;
      RECT 1139.000000 660.350000 1149.500000 663.650000 ;
      RECT 657.500000 660.350000 658.500000 661.650000 ;
      RECT 616.500000 660.350000 649.500000 661.650000 ;
      RECT 607.500000 660.350000 608.500000 661.650000 ;
      RECT 566.500000 660.350000 599.500000 661.650000 ;
      RECT 557.500000 660.350000 558.500000 661.650000 ;
      RECT 516.500000 660.350000 549.500000 661.650000 ;
      RECT 507.500000 660.350000 508.500000 661.650000 ;
      RECT 466.500000 660.350000 499.500000 661.650000 ;
      RECT 457.500000 660.350000 458.500000 661.650000 ;
      RECT 416.500000 660.350000 449.500000 661.650000 ;
      RECT 407.500000 660.350000 408.500000 661.650000 ;
      RECT 396.500000 660.350000 399.500000 663.650000 ;
      RECT 382.500000 660.350000 383.500000 661.650000 ;
      RECT 357.500000 660.350000 358.500000 661.650000 ;
      RECT 2.020000 660.350000 349.500000 663.170000 ;
      RECT 2.020000 660.070000 358.500000 660.350000 ;
      RECT 1166.500000 660.065000 1183.980000 661.650000 ;
      RECT 1139.000000 659.650000 1158.500000 660.350000 ;
      RECT 616.500000 659.650000 658.500000 660.350000 ;
      RECT 566.500000 659.650000 608.500000 660.350000 ;
      RECT 516.500000 659.650000 558.500000 660.350000 ;
      RECT 466.500000 659.650000 508.500000 660.350000 ;
      RECT 416.500000 659.650000 458.500000 660.350000 ;
      RECT 382.500000 659.650000 408.500000 660.350000 ;
      RECT 0.000000 659.650000 358.500000 660.070000 ;
      RECT 1166.500000 658.350000 1186.000000 660.065000 ;
      RECT 1157.500000 658.350000 1158.500000 659.650000 ;
      RECT 666.500000 658.350000 670.000000 661.650000 ;
      RECT 657.500000 658.350000 658.500000 659.650000 ;
      RECT 616.500000 658.350000 649.500000 659.650000 ;
      RECT 607.500000 658.350000 608.500000 659.650000 ;
      RECT 566.500000 658.350000 599.500000 659.650000 ;
      RECT 557.500000 658.350000 558.500000 659.650000 ;
      RECT 516.500000 658.350000 549.500000 659.650000 ;
      RECT 507.500000 658.350000 508.500000 659.650000 ;
      RECT 466.500000 658.350000 499.500000 659.650000 ;
      RECT 457.500000 658.350000 458.500000 659.650000 ;
      RECT 416.500000 658.350000 449.500000 659.650000 ;
      RECT 407.500000 658.350000 408.500000 659.650000 ;
      RECT 382.500000 658.350000 383.500000 659.650000 ;
      RECT 366.500000 658.350000 369.500000 661.650000 ;
      RECT 357.500000 658.350000 358.500000 659.650000 ;
      RECT 1157.500000 657.650000 1186.000000 658.350000 ;
      RECT 357.500000 657.650000 383.500000 658.350000 ;
      RECT 1166.500000 657.485000 1186.000000 657.650000 ;
      RECT 1157.500000 656.350000 1158.500000 657.650000 ;
      RECT 1139.000000 656.350000 1149.500000 659.650000 ;
      RECT 657.500000 656.350000 670.000000 658.350000 ;
      RECT 607.500000 656.350000 649.500000 658.350000 ;
      RECT 557.500000 656.350000 599.500000 658.350000 ;
      RECT 507.500000 656.350000 549.500000 658.350000 ;
      RECT 457.500000 656.350000 499.500000 658.350000 ;
      RECT 407.500000 656.350000 449.500000 658.350000 ;
      RECT 396.500000 656.350000 399.500000 659.650000 ;
      RECT 382.500000 656.350000 383.500000 657.650000 ;
      RECT 357.500000 656.350000 358.500000 657.650000 ;
      RECT 0.000000 656.350000 349.500000 659.650000 ;
      RECT 382.500000 656.000000 670.000000 656.350000 ;
      RECT 1139.000000 655.650000 1158.500000 656.350000 ;
      RECT 382.500000 655.650000 399.000000 656.000000 ;
      RECT 0.000000 655.650000 358.500000 656.350000 ;
      RECT 1166.500000 654.385000 1183.980000 657.485000 ;
      RECT 1166.500000 654.350000 1186.000000 654.385000 ;
      RECT 1157.500000 654.350000 1158.500000 655.650000 ;
      RECT 382.500000 654.350000 383.500000 655.650000 ;
      RECT 366.500000 654.350000 369.500000 657.650000 ;
      RECT 357.500000 654.350000 358.500000 655.650000 ;
      RECT 1157.500000 653.650000 1186.000000 654.350000 ;
      RECT 357.500000 653.650000 383.500000 654.350000 ;
      RECT 1166.500000 653.525000 1186.000000 653.650000 ;
      RECT 0.000000 652.575000 349.500000 655.650000 ;
      RECT 1157.500000 652.350000 1158.500000 653.650000 ;
      RECT 1139.000000 652.350000 1149.500000 655.650000 ;
      RECT 396.500000 652.350000 399.000000 655.650000 ;
      RECT 382.500000 652.350000 383.500000 653.650000 ;
      RECT 357.500000 652.350000 358.500000 653.650000 ;
      RECT 2.020000 652.350000 349.500000 652.575000 ;
      RECT 1139.000000 651.650000 1158.500000 652.350000 ;
      RECT 382.500000 651.650000 399.000000 652.350000 ;
      RECT 2.020000 651.650000 358.500000 652.350000 ;
      RECT 1166.500000 650.425000 1183.980000 653.525000 ;
      RECT 1166.500000 650.350000 1186.000000 650.425000 ;
      RECT 1157.500000 650.350000 1158.500000 651.650000 ;
      RECT 382.500000 650.350000 383.500000 651.650000 ;
      RECT 366.500000 650.350000 369.500000 653.650000 ;
      RECT 357.500000 650.350000 358.500000 651.650000 ;
      RECT 1157.500000 649.650000 1186.000000 650.350000 ;
      RECT 357.500000 649.650000 383.500000 650.350000 ;
      RECT 2.020000 649.475000 349.500000 651.650000 ;
      RECT 0.000000 648.615000 349.500000 649.475000 ;
      RECT 1157.500000 648.350000 1158.500000 649.650000 ;
      RECT 1139.000000 648.350000 1149.500000 651.650000 ;
      RECT 396.500000 648.350000 399.000000 651.650000 ;
      RECT 382.500000 648.350000 383.500000 649.650000 ;
      RECT 357.500000 648.350000 358.500000 649.650000 ;
      RECT 2.020000 648.350000 349.500000 648.615000 ;
      RECT 1139.000000 647.650000 1158.500000 648.350000 ;
      RECT 382.500000 647.650000 399.000000 648.350000 ;
      RECT 2.020000 647.650000 358.500000 648.350000 ;
      RECT 1166.500000 646.350000 1186.000000 649.650000 ;
      RECT 1157.500000 646.350000 1158.500000 647.650000 ;
      RECT 382.500000 646.350000 383.500000 647.650000 ;
      RECT 366.500000 646.350000 369.500000 649.650000 ;
      RECT 357.500000 646.350000 358.500000 647.650000 ;
      RECT 1157.500000 645.650000 1186.000000 646.350000 ;
      RECT 357.500000 645.650000 383.500000 646.350000 ;
      RECT 2.020000 645.515000 349.500000 647.650000 ;
      RECT 1157.500000 644.350000 1158.500000 645.650000 ;
      RECT 1139.000000 644.350000 1149.500000 647.650000 ;
      RECT 396.500000 644.350000 399.000000 647.650000 ;
      RECT 382.500000 644.350000 383.500000 645.650000 ;
      RECT 357.500000 644.350000 358.500000 645.650000 ;
      RECT 0.000000 644.350000 349.500000 645.515000 ;
      RECT 1139.000000 643.650000 1158.500000 644.350000 ;
      RECT 382.500000 643.650000 399.000000 644.350000 ;
      RECT 0.000000 643.650000 358.500000 644.350000 ;
      RECT 0.000000 642.935000 349.500000 643.650000 ;
      RECT 1166.500000 642.930000 1186.000000 645.650000 ;
      RECT 1166.500000 642.350000 1183.980000 642.930000 ;
      RECT 1157.500000 642.350000 1158.500000 643.650000 ;
      RECT 382.500000 642.350000 383.500000 643.650000 ;
      RECT 366.500000 642.350000 369.500000 645.650000 ;
      RECT 357.500000 642.350000 358.500000 643.650000 ;
      RECT 1157.500000 641.650000 1183.980000 642.350000 ;
      RECT 357.500000 641.650000 383.500000 642.350000 ;
      RECT 1157.500000 640.350000 1158.500000 641.650000 ;
      RECT 1139.000000 640.350000 1149.500000 643.650000 ;
      RECT 396.500000 640.350000 399.000000 643.650000 ;
      RECT 382.500000 640.350000 383.500000 641.650000 ;
      RECT 357.500000 640.350000 358.500000 641.650000 ;
      RECT 2.020000 640.350000 349.500000 642.935000 ;
      RECT 2.020000 639.835000 358.500000 640.350000 ;
      RECT 1166.500000 639.830000 1183.980000 641.650000 ;
      RECT 1139.000000 639.650000 1158.500000 640.350000 ;
      RECT 382.500000 639.650000 399.000000 640.350000 ;
      RECT 0.000000 639.650000 358.500000 639.835000 ;
      RECT 1166.500000 638.350000 1186.000000 639.830000 ;
      RECT 1157.500000 638.350000 1158.500000 639.650000 ;
      RECT 382.500000 638.350000 383.500000 639.650000 ;
      RECT 366.500000 638.350000 369.500000 641.650000 ;
      RECT 357.500000 638.350000 358.500000 639.650000 ;
      RECT 1157.500000 637.650000 1186.000000 638.350000 ;
      RECT 357.500000 637.650000 383.500000 638.350000 ;
      RECT 1157.500000 636.350000 1158.500000 637.650000 ;
      RECT 1139.000000 636.350000 1149.500000 639.650000 ;
      RECT 396.500000 636.350000 399.000000 639.650000 ;
      RECT 382.500000 636.350000 383.500000 637.650000 ;
      RECT 357.500000 636.350000 358.500000 637.650000 ;
      RECT 0.000000 636.350000 349.500000 639.650000 ;
      RECT 1139.000000 635.650000 1158.500000 636.350000 ;
      RECT 382.500000 635.650000 399.000000 636.350000 ;
      RECT 0.000000 635.650000 358.500000 636.350000 ;
      RECT 1166.500000 634.350000 1186.000000 637.650000 ;
      RECT 1157.500000 634.350000 1158.500000 635.650000 ;
      RECT 382.500000 634.350000 383.500000 635.650000 ;
      RECT 366.500000 634.350000 369.500000 637.650000 ;
      RECT 357.500000 634.350000 358.500000 635.650000 ;
      RECT 1157.500000 633.650000 1186.000000 634.350000 ;
      RECT 357.500000 633.650000 383.500000 634.350000 ;
      RECT 1157.500000 632.350000 1158.500000 633.650000 ;
      RECT 1139.000000 632.350000 1149.500000 635.650000 ;
      RECT 396.500000 632.350000 399.000000 635.650000 ;
      RECT 382.500000 632.350000 383.500000 633.650000 ;
      RECT 357.500000 632.350000 358.500000 633.650000 ;
      RECT 0.000000 632.350000 349.500000 635.650000 ;
      RECT 1139.000000 631.650000 1158.500000 632.350000 ;
      RECT 382.500000 631.650000 399.000000 632.350000 ;
      RECT 0.000000 631.650000 358.500000 632.350000 ;
      RECT 1166.500000 630.350000 1186.000000 633.650000 ;
      RECT 1157.500000 630.350000 1158.500000 631.650000 ;
      RECT 382.500000 630.350000 383.500000 631.650000 ;
      RECT 366.500000 630.350000 369.500000 633.650000 ;
      RECT 357.500000 630.350000 358.500000 631.650000 ;
      RECT 1157.500000 629.650000 1186.000000 630.350000 ;
      RECT 357.500000 629.650000 383.500000 630.350000 ;
      RECT 1157.500000 628.350000 1158.500000 629.650000 ;
      RECT 1139.000000 628.350000 1149.500000 631.650000 ;
      RECT 396.500000 628.350000 399.000000 631.650000 ;
      RECT 382.500000 628.350000 383.500000 629.650000 ;
      RECT 357.500000 628.350000 358.500000 629.650000 ;
      RECT 0.000000 628.350000 349.500000 631.650000 ;
      RECT 1139.000000 627.650000 1158.500000 628.350000 ;
      RECT 382.500000 627.650000 399.000000 628.350000 ;
      RECT 0.000000 627.650000 358.500000 628.350000 ;
      RECT 1166.500000 626.350000 1186.000000 629.650000 ;
      RECT 1157.500000 626.350000 1158.500000 627.650000 ;
      RECT 382.500000 626.350000 383.500000 627.650000 ;
      RECT 366.500000 626.350000 369.500000 629.650000 ;
      RECT 357.500000 626.350000 358.500000 627.650000 ;
      RECT 1157.500000 625.650000 1186.000000 626.350000 ;
      RECT 357.500000 625.650000 383.500000 626.350000 ;
      RECT 1157.500000 624.350000 1158.500000 625.650000 ;
      RECT 1139.000000 624.350000 1149.500000 627.650000 ;
      RECT 396.500000 624.350000 399.000000 627.650000 ;
      RECT 382.500000 624.350000 383.500000 625.650000 ;
      RECT 357.500000 624.350000 358.500000 625.650000 ;
      RECT 0.000000 624.350000 349.500000 627.650000 ;
      RECT 1139.000000 623.650000 1158.500000 624.350000 ;
      RECT 382.500000 623.650000 399.000000 624.350000 ;
      RECT 0.000000 623.650000 358.500000 624.350000 ;
      RECT 1166.500000 622.350000 1186.000000 625.650000 ;
      RECT 1157.500000 622.350000 1158.500000 623.650000 ;
      RECT 382.500000 622.350000 383.500000 623.650000 ;
      RECT 366.500000 622.350000 369.500000 625.650000 ;
      RECT 357.500000 622.350000 358.500000 623.650000 ;
      RECT 1157.500000 621.650000 1186.000000 622.350000 ;
      RECT 357.500000 621.650000 383.500000 622.350000 ;
      RECT 1157.500000 620.350000 1158.500000 621.650000 ;
      RECT 1139.000000 620.350000 1149.500000 623.650000 ;
      RECT 396.500000 620.350000 399.000000 623.650000 ;
      RECT 382.500000 620.350000 383.500000 621.650000 ;
      RECT 357.500000 620.350000 358.500000 621.650000 ;
      RECT 0.000000 620.350000 349.500000 623.650000 ;
      RECT 1139.000000 619.650000 1158.500000 620.350000 ;
      RECT 382.500000 619.650000 399.000000 620.350000 ;
      RECT 0.000000 619.650000 358.500000 620.350000 ;
      RECT 1166.500000 618.350000 1186.000000 621.650000 ;
      RECT 1157.500000 618.350000 1158.500000 619.650000 ;
      RECT 382.500000 618.350000 383.500000 619.650000 ;
      RECT 366.500000 618.350000 369.500000 621.650000 ;
      RECT 357.500000 618.350000 358.500000 619.650000 ;
      RECT 1157.500000 617.650000 1186.000000 618.350000 ;
      RECT 357.500000 617.650000 383.500000 618.350000 ;
      RECT 1157.500000 616.350000 1158.500000 617.650000 ;
      RECT 1139.000000 616.350000 1149.500000 619.650000 ;
      RECT 396.500000 616.350000 399.000000 619.650000 ;
      RECT 382.500000 616.350000 383.500000 617.650000 ;
      RECT 357.500000 616.350000 358.500000 617.650000 ;
      RECT 0.000000 616.350000 349.500000 619.650000 ;
      RECT 382.500000 616.115000 399.000000 616.350000 ;
      RECT 1139.000000 615.695000 1158.500000 616.350000 ;
      RECT 1141.020000 615.650000 1158.500000 615.695000 ;
      RECT 382.500000 615.650000 396.980000 616.115000 ;
      RECT 0.000000 615.650000 358.500000 616.350000 ;
      RECT 1166.500000 614.350000 1186.000000 617.650000 ;
      RECT 1157.500000 614.350000 1158.500000 615.650000 ;
      RECT 382.500000 614.350000 383.500000 615.650000 ;
      RECT 366.500000 614.350000 369.500000 617.650000 ;
      RECT 357.500000 614.350000 358.500000 615.650000 ;
      RECT 1157.500000 613.650000 1186.000000 614.350000 ;
      RECT 357.500000 613.650000 383.500000 614.350000 ;
      RECT 1157.500000 612.350000 1158.500000 613.650000 ;
      RECT 1141.020000 612.350000 1149.500000 615.650000 ;
      RECT 396.500000 612.350000 396.980000 615.650000 ;
      RECT 382.500000 612.350000 383.500000 613.650000 ;
      RECT 357.500000 612.350000 358.500000 613.650000 ;
      RECT 0.000000 612.350000 349.500000 615.650000 ;
      RECT 1141.020000 611.650000 1158.500000 612.350000 ;
      RECT 382.500000 611.650000 396.980000 612.350000 ;
      RECT 0.000000 611.650000 358.500000 612.350000 ;
      RECT 1166.500000 610.350000 1186.000000 613.650000 ;
      RECT 1157.500000 610.350000 1158.500000 611.650000 ;
      RECT 382.500000 610.350000 383.500000 611.650000 ;
      RECT 366.500000 610.350000 369.500000 613.650000 ;
      RECT 357.500000 610.350000 358.500000 611.650000 ;
      RECT 1157.500000 609.650000 1186.000000 610.350000 ;
      RECT 357.500000 609.650000 383.500000 610.350000 ;
      RECT 1157.500000 608.350000 1158.500000 609.650000 ;
      RECT 1141.020000 608.350000 1149.500000 611.650000 ;
      RECT 396.500000 608.350000 396.980000 611.650000 ;
      RECT 382.500000 608.350000 383.500000 609.650000 ;
      RECT 357.500000 608.350000 358.500000 609.650000 ;
      RECT 0.000000 608.350000 349.500000 611.650000 ;
      RECT 1141.020000 607.650000 1158.500000 608.350000 ;
      RECT 382.500000 607.650000 396.980000 608.350000 ;
      RECT 0.000000 607.650000 358.500000 608.350000 ;
      RECT 1166.500000 606.350000 1186.000000 609.650000 ;
      RECT 1157.500000 606.350000 1158.500000 607.650000 ;
      RECT 382.500000 606.350000 383.500000 607.650000 ;
      RECT 366.500000 606.350000 369.500000 609.650000 ;
      RECT 357.500000 606.350000 358.500000 607.650000 ;
      RECT 1157.500000 605.650000 1186.000000 606.350000 ;
      RECT 357.500000 605.650000 383.500000 606.350000 ;
      RECT 1157.500000 604.350000 1158.500000 605.650000 ;
      RECT 1141.020000 604.350000 1149.500000 607.650000 ;
      RECT 396.500000 604.350000 396.980000 607.650000 ;
      RECT 382.500000 604.350000 383.500000 605.650000 ;
      RECT 357.500000 604.350000 358.500000 605.650000 ;
      RECT 0.000000 604.350000 349.500000 607.650000 ;
      RECT 1141.020000 603.650000 1158.500000 604.350000 ;
      RECT 382.500000 603.650000 396.980000 604.350000 ;
      RECT 0.000000 603.650000 358.500000 604.350000 ;
      RECT 1166.500000 602.350000 1186.000000 605.650000 ;
      RECT 1157.500000 602.350000 1158.500000 603.650000 ;
      RECT 382.500000 602.350000 383.500000 603.650000 ;
      RECT 366.500000 602.350000 369.500000 605.650000 ;
      RECT 357.500000 602.350000 358.500000 603.650000 ;
      RECT 1157.500000 601.650000 1186.000000 602.350000 ;
      RECT 357.500000 601.650000 383.500000 602.350000 ;
      RECT 1157.500000 600.350000 1158.500000 601.650000 ;
      RECT 1141.020000 600.350000 1149.500000 603.650000 ;
      RECT 396.500000 600.350000 396.980000 603.650000 ;
      RECT 382.500000 600.350000 383.500000 601.650000 ;
      RECT 357.500000 600.350000 358.500000 601.650000 ;
      RECT 0.000000 600.350000 349.500000 603.650000 ;
      RECT 1141.020000 599.650000 1158.500000 600.350000 ;
      RECT 382.500000 599.650000 396.980000 600.350000 ;
      RECT 0.000000 599.650000 358.500000 600.350000 ;
      RECT 1166.500000 598.350000 1186.000000 601.650000 ;
      RECT 1157.500000 598.350000 1158.500000 599.650000 ;
      RECT 382.500000 598.350000 383.500000 599.650000 ;
      RECT 366.500000 598.350000 369.500000 601.650000 ;
      RECT 357.500000 598.350000 358.500000 599.650000 ;
      RECT 1141.020000 597.880000 1149.500000 599.650000 ;
      RECT 1157.500000 597.650000 1186.000000 598.350000 ;
      RECT 357.500000 597.650000 383.500000 598.350000 ;
      RECT 1157.500000 596.350000 1158.500000 597.650000 ;
      RECT 1139.000000 596.350000 1149.500000 597.880000 ;
      RECT 396.500000 596.350000 396.980000 599.650000 ;
      RECT 382.500000 596.350000 383.500000 597.650000 ;
      RECT 357.500000 596.350000 358.500000 597.650000 ;
      RECT 0.000000 596.350000 349.500000 599.650000 ;
      RECT 1139.000000 595.650000 1158.500000 596.350000 ;
      RECT 382.500000 595.650000 396.980000 596.350000 ;
      RECT 0.000000 595.650000 358.500000 596.350000 ;
      RECT 1166.500000 594.350000 1186.000000 597.650000 ;
      RECT 1157.500000 594.350000 1158.500000 595.650000 ;
      RECT 382.500000 594.350000 383.500000 595.650000 ;
      RECT 366.500000 594.350000 369.500000 597.650000 ;
      RECT 357.500000 594.350000 358.500000 595.650000 ;
      RECT 1157.500000 593.650000 1186.000000 594.350000 ;
      RECT 357.500000 593.650000 383.500000 594.350000 ;
      RECT 1157.500000 592.350000 1158.500000 593.650000 ;
      RECT 1139.000000 592.350000 1149.500000 595.650000 ;
      RECT 396.500000 592.350000 396.980000 595.650000 ;
      RECT 382.500000 592.350000 383.500000 593.650000 ;
      RECT 357.500000 592.350000 358.500000 593.650000 ;
      RECT 0.000000 592.350000 349.500000 595.650000 ;
      RECT 1139.000000 591.650000 1158.500000 592.350000 ;
      RECT 382.500000 591.650000 396.980000 592.350000 ;
      RECT 0.000000 591.650000 358.500000 592.350000 ;
      RECT 1166.500000 590.350000 1186.000000 593.650000 ;
      RECT 1157.500000 590.350000 1158.500000 591.650000 ;
      RECT 382.500000 590.350000 383.500000 591.650000 ;
      RECT 366.500000 590.350000 369.500000 593.650000 ;
      RECT 357.500000 590.350000 358.500000 591.650000 ;
      RECT 1157.500000 589.650000 1186.000000 590.350000 ;
      RECT 357.500000 589.650000 383.500000 590.350000 ;
      RECT 1157.500000 588.350000 1158.500000 589.650000 ;
      RECT 1139.000000 588.350000 1149.500000 591.650000 ;
      RECT 396.500000 588.350000 396.980000 591.650000 ;
      RECT 382.500000 588.350000 383.500000 589.650000 ;
      RECT 357.500000 588.350000 358.500000 589.650000 ;
      RECT 0.000000 588.350000 349.500000 591.650000 ;
      RECT 1139.000000 587.650000 1158.500000 588.350000 ;
      RECT 382.500000 587.650000 396.980000 588.350000 ;
      RECT 0.000000 587.650000 358.500000 588.350000 ;
      RECT 1166.500000 586.350000 1186.000000 589.650000 ;
      RECT 1157.500000 586.350000 1158.500000 587.650000 ;
      RECT 382.500000 586.350000 383.500000 587.650000 ;
      RECT 366.500000 586.350000 369.500000 589.650000 ;
      RECT 357.500000 586.350000 358.500000 587.650000 ;
      RECT 1157.500000 585.650000 1186.000000 586.350000 ;
      RECT 357.500000 585.650000 383.500000 586.350000 ;
      RECT 1157.500000 584.350000 1158.500000 585.650000 ;
      RECT 1139.000000 584.350000 1149.500000 587.650000 ;
      RECT 396.500000 584.350000 396.980000 587.650000 ;
      RECT 382.500000 584.350000 383.500000 585.650000 ;
      RECT 357.500000 584.350000 358.500000 585.650000 ;
      RECT 0.000000 584.350000 349.500000 587.650000 ;
      RECT 1139.000000 583.650000 1158.500000 584.350000 ;
      RECT 382.500000 583.650000 396.980000 584.350000 ;
      RECT 0.000000 583.650000 358.500000 584.350000 ;
      RECT 1166.500000 582.350000 1186.000000 585.650000 ;
      RECT 1157.500000 582.350000 1158.500000 583.650000 ;
      RECT 382.500000 582.350000 383.500000 583.650000 ;
      RECT 366.500000 582.350000 369.500000 585.650000 ;
      RECT 357.500000 582.350000 358.500000 583.650000 ;
      RECT 1157.500000 581.650000 1186.000000 582.350000 ;
      RECT 357.500000 581.650000 383.500000 582.350000 ;
      RECT 1157.500000 580.350000 1158.500000 581.650000 ;
      RECT 1139.000000 580.350000 1149.500000 583.650000 ;
      RECT 396.500000 580.350000 396.980000 583.650000 ;
      RECT 382.500000 580.350000 383.500000 581.650000 ;
      RECT 357.500000 580.350000 358.500000 581.650000 ;
      RECT 0.000000 580.350000 349.500000 583.650000 ;
      RECT 1139.000000 579.650000 1158.500000 580.350000 ;
      RECT 382.500000 579.650000 396.980000 580.350000 ;
      RECT 0.000000 579.650000 358.500000 580.350000 ;
      RECT 1166.500000 578.350000 1186.000000 581.650000 ;
      RECT 1157.500000 578.350000 1158.500000 579.650000 ;
      RECT 382.500000 578.350000 383.500000 579.650000 ;
      RECT 366.500000 578.350000 369.500000 581.650000 ;
      RECT 357.500000 578.350000 358.500000 579.650000 ;
      RECT 1157.500000 577.650000 1186.000000 578.350000 ;
      RECT 357.500000 577.650000 383.500000 578.350000 ;
      RECT 396.500000 577.590000 396.980000 579.650000 ;
      RECT 1157.500000 576.350000 1158.500000 577.650000 ;
      RECT 1139.000000 576.350000 1149.500000 579.650000 ;
      RECT 396.500000 576.350000 399.000000 577.590000 ;
      RECT 382.500000 576.350000 383.500000 577.650000 ;
      RECT 357.500000 576.350000 358.500000 577.650000 ;
      RECT 0.000000 576.350000 349.500000 579.650000 ;
      RECT 1139.000000 575.650000 1158.500000 576.350000 ;
      RECT 382.500000 575.650000 399.000000 576.350000 ;
      RECT 0.000000 575.650000 358.500000 576.350000 ;
      RECT 0.000000 575.170000 349.500000 575.650000 ;
      RECT 1166.500000 575.165000 1186.000000 577.650000 ;
      RECT 1166.500000 574.350000 1183.980000 575.165000 ;
      RECT 1157.500000 574.350000 1158.500000 575.650000 ;
      RECT 382.500000 574.350000 383.500000 575.650000 ;
      RECT 366.500000 574.350000 369.500000 577.650000 ;
      RECT 357.500000 574.350000 358.500000 575.650000 ;
      RECT 1157.500000 573.650000 1183.980000 574.350000 ;
      RECT 357.500000 573.650000 383.500000 574.350000 ;
      RECT 1157.500000 572.350000 1158.500000 573.650000 ;
      RECT 1139.000000 572.350000 1149.500000 575.650000 ;
      RECT 396.500000 572.350000 399.000000 575.650000 ;
      RECT 382.500000 572.350000 383.500000 573.650000 ;
      RECT 357.500000 572.350000 358.500000 573.650000 ;
      RECT 2.020000 572.350000 349.500000 575.170000 ;
      RECT 2.020000 572.070000 358.500000 572.350000 ;
      RECT 1166.500000 572.065000 1183.980000 573.650000 ;
      RECT 1139.000000 571.650000 1158.500000 572.350000 ;
      RECT 382.500000 571.650000 399.000000 572.350000 ;
      RECT 0.000000 571.650000 358.500000 572.070000 ;
      RECT 1166.500000 570.350000 1186.000000 572.065000 ;
      RECT 1157.500000 570.350000 1158.500000 571.650000 ;
      RECT 382.500000 570.350000 383.500000 571.650000 ;
      RECT 366.500000 570.350000 369.500000 573.650000 ;
      RECT 357.500000 570.350000 358.500000 571.650000 ;
      RECT 1157.500000 569.650000 1186.000000 570.350000 ;
      RECT 357.500000 569.650000 383.500000 570.350000 ;
      RECT 1166.500000 569.485000 1186.000000 569.650000 ;
      RECT 1157.500000 568.350000 1158.500000 569.650000 ;
      RECT 1139.000000 568.350000 1149.500000 571.650000 ;
      RECT 396.500000 568.350000 399.000000 571.650000 ;
      RECT 382.500000 568.350000 383.500000 569.650000 ;
      RECT 357.500000 568.350000 358.500000 569.650000 ;
      RECT 0.000000 568.350000 349.500000 571.650000 ;
      RECT 1139.000000 567.650000 1158.500000 568.350000 ;
      RECT 382.500000 567.650000 399.000000 568.350000 ;
      RECT 0.000000 567.650000 358.500000 568.350000 ;
      RECT 1166.500000 566.385000 1183.980000 569.485000 ;
      RECT 1166.500000 566.350000 1186.000000 566.385000 ;
      RECT 1157.500000 566.350000 1158.500000 567.650000 ;
      RECT 382.500000 566.350000 383.500000 567.650000 ;
      RECT 366.500000 566.350000 369.500000 569.650000 ;
      RECT 357.500000 566.350000 358.500000 567.650000 ;
      RECT 1157.500000 565.650000 1186.000000 566.350000 ;
      RECT 357.500000 565.650000 383.500000 566.350000 ;
      RECT 1166.500000 565.525000 1186.000000 565.650000 ;
      RECT 0.000000 564.575000 349.500000 567.650000 ;
      RECT 1157.500000 564.350000 1158.500000 565.650000 ;
      RECT 1139.000000 564.350000 1149.500000 567.650000 ;
      RECT 396.500000 564.350000 399.000000 567.650000 ;
      RECT 382.500000 564.350000 383.500000 565.650000 ;
      RECT 357.500000 564.350000 358.500000 565.650000 ;
      RECT 2.020000 564.350000 349.500000 564.575000 ;
      RECT 1139.000000 563.650000 1158.500000 564.350000 ;
      RECT 382.500000 563.650000 399.000000 564.350000 ;
      RECT 2.020000 563.650000 358.500000 564.350000 ;
      RECT 1166.500000 562.425000 1183.980000 565.525000 ;
      RECT 1166.500000 562.350000 1186.000000 562.425000 ;
      RECT 1157.500000 562.350000 1158.500000 563.650000 ;
      RECT 382.500000 562.350000 383.500000 563.650000 ;
      RECT 366.500000 562.350000 369.500000 565.650000 ;
      RECT 357.500000 562.350000 358.500000 563.650000 ;
      RECT 1157.500000 561.650000 1186.000000 562.350000 ;
      RECT 357.500000 561.650000 383.500000 562.350000 ;
      RECT 2.020000 561.475000 349.500000 563.650000 ;
      RECT 0.000000 560.615000 349.500000 561.475000 ;
      RECT 1157.500000 560.350000 1158.500000 561.650000 ;
      RECT 1139.000000 560.350000 1149.500000 563.650000 ;
      RECT 396.500000 560.350000 399.000000 563.650000 ;
      RECT 382.500000 560.350000 383.500000 561.650000 ;
      RECT 357.500000 560.350000 358.500000 561.650000 ;
      RECT 2.020000 560.350000 349.500000 560.615000 ;
      RECT 1139.000000 559.650000 1158.500000 560.350000 ;
      RECT 382.500000 559.650000 399.000000 560.350000 ;
      RECT 2.020000 559.650000 358.500000 560.350000 ;
      RECT 1166.500000 558.350000 1186.000000 561.650000 ;
      RECT 1157.500000 558.350000 1158.500000 559.650000 ;
      RECT 382.500000 558.350000 383.500000 559.650000 ;
      RECT 366.500000 558.350000 369.500000 561.650000 ;
      RECT 357.500000 558.350000 358.500000 559.650000 ;
      RECT 1157.500000 557.650000 1186.000000 558.350000 ;
      RECT 357.500000 557.650000 383.500000 558.350000 ;
      RECT 2.020000 557.515000 349.500000 559.650000 ;
      RECT 1157.500000 556.350000 1158.500000 557.650000 ;
      RECT 1139.000000 556.350000 1149.500000 559.650000 ;
      RECT 396.500000 556.350000 399.000000 559.650000 ;
      RECT 382.500000 556.350000 383.500000 557.650000 ;
      RECT 357.500000 556.350000 358.500000 557.650000 ;
      RECT 0.000000 556.350000 349.500000 557.515000 ;
      RECT 1139.000000 555.650000 1158.500000 556.350000 ;
      RECT 382.500000 555.650000 399.000000 556.350000 ;
      RECT 0.000000 555.650000 358.500000 556.350000 ;
      RECT 0.000000 554.935000 349.500000 555.650000 ;
      RECT 1166.500000 554.930000 1186.000000 557.650000 ;
      RECT 1166.500000 554.350000 1183.980000 554.930000 ;
      RECT 1157.500000 554.350000 1158.500000 555.650000 ;
      RECT 382.500000 554.350000 383.500000 555.650000 ;
      RECT 366.500000 554.350000 369.500000 557.650000 ;
      RECT 357.500000 554.350000 358.500000 555.650000 ;
      RECT 1157.500000 553.650000 1183.980000 554.350000 ;
      RECT 357.500000 553.650000 383.500000 554.350000 ;
      RECT 1157.500000 552.350000 1158.500000 553.650000 ;
      RECT 1139.000000 552.350000 1149.500000 555.650000 ;
      RECT 396.500000 552.350000 399.000000 555.650000 ;
      RECT 382.500000 552.350000 383.500000 553.650000 ;
      RECT 357.500000 552.350000 358.500000 553.650000 ;
      RECT 2.020000 552.350000 349.500000 554.935000 ;
      RECT 2.020000 551.835000 358.500000 552.350000 ;
      RECT 1166.500000 551.830000 1183.980000 553.650000 ;
      RECT 1139.000000 551.650000 1158.500000 552.350000 ;
      RECT 382.500000 551.650000 399.000000 552.350000 ;
      RECT 0.000000 551.650000 358.500000 551.835000 ;
      RECT 1166.500000 550.350000 1186.000000 551.830000 ;
      RECT 1157.500000 550.350000 1158.500000 551.650000 ;
      RECT 382.500000 550.350000 383.500000 551.650000 ;
      RECT 366.500000 550.350000 369.500000 553.650000 ;
      RECT 357.500000 550.350000 358.500000 551.650000 ;
      RECT 1157.500000 549.650000 1186.000000 550.350000 ;
      RECT 357.500000 549.650000 383.500000 550.350000 ;
      RECT 1157.500000 548.350000 1158.500000 549.650000 ;
      RECT 1139.000000 548.350000 1149.500000 551.650000 ;
      RECT 396.500000 548.350000 399.000000 551.650000 ;
      RECT 382.500000 548.350000 383.500000 549.650000 ;
      RECT 357.500000 548.350000 358.500000 549.650000 ;
      RECT 0.000000 548.350000 349.500000 551.650000 ;
      RECT 1139.000000 547.650000 1158.500000 548.350000 ;
      RECT 382.500000 547.650000 399.000000 548.350000 ;
      RECT 0.000000 547.650000 358.500000 548.350000 ;
      RECT 1166.500000 546.350000 1186.000000 549.650000 ;
      RECT 1157.500000 546.350000 1158.500000 547.650000 ;
      RECT 382.500000 546.350000 383.500000 547.650000 ;
      RECT 366.500000 546.350000 369.500000 549.650000 ;
      RECT 357.500000 546.350000 358.500000 547.650000 ;
      RECT 1157.500000 545.650000 1186.000000 546.350000 ;
      RECT 357.500000 545.650000 383.500000 546.350000 ;
      RECT 1157.500000 544.350000 1158.500000 545.650000 ;
      RECT 1139.000000 544.350000 1149.500000 547.650000 ;
      RECT 396.500000 544.350000 399.000000 547.650000 ;
      RECT 382.500000 544.350000 383.500000 545.650000 ;
      RECT 357.500000 544.350000 358.500000 545.650000 ;
      RECT 0.000000 544.350000 349.500000 547.650000 ;
      RECT 1139.000000 543.650000 1158.500000 544.350000 ;
      RECT 382.500000 543.650000 399.000000 544.350000 ;
      RECT 0.000000 543.650000 358.500000 544.350000 ;
      RECT 1166.500000 542.350000 1186.000000 545.650000 ;
      RECT 1157.500000 542.350000 1158.500000 543.650000 ;
      RECT 382.500000 542.350000 383.500000 543.650000 ;
      RECT 366.500000 542.350000 369.500000 545.650000 ;
      RECT 357.500000 542.350000 358.500000 543.650000 ;
      RECT 1157.500000 541.650000 1186.000000 542.350000 ;
      RECT 357.500000 541.650000 383.500000 542.350000 ;
      RECT 1157.500000 540.350000 1158.500000 541.650000 ;
      RECT 1139.000000 540.350000 1149.500000 543.650000 ;
      RECT 396.500000 540.350000 399.000000 543.650000 ;
      RECT 382.500000 540.350000 383.500000 541.650000 ;
      RECT 357.500000 540.350000 358.500000 541.650000 ;
      RECT 0.000000 540.350000 349.500000 543.650000 ;
      RECT 1139.000000 539.650000 1158.500000 540.350000 ;
      RECT 382.500000 539.650000 399.000000 540.350000 ;
      RECT 0.000000 539.650000 358.500000 540.350000 ;
      RECT 1166.500000 538.350000 1186.000000 541.650000 ;
      RECT 1157.500000 538.350000 1158.500000 539.650000 ;
      RECT 382.500000 538.350000 383.500000 539.650000 ;
      RECT 366.500000 538.350000 369.500000 541.650000 ;
      RECT 357.500000 538.350000 358.500000 539.650000 ;
      RECT 1157.500000 537.650000 1186.000000 538.350000 ;
      RECT 357.500000 537.650000 383.500000 538.350000 ;
      RECT 1157.500000 536.350000 1158.500000 537.650000 ;
      RECT 1139.000000 536.350000 1149.500000 539.650000 ;
      RECT 396.500000 536.350000 399.000000 539.650000 ;
      RECT 382.500000 536.350000 383.500000 537.650000 ;
      RECT 357.500000 536.350000 358.500000 537.650000 ;
      RECT 0.000000 536.350000 349.500000 539.650000 ;
      RECT 1139.000000 535.650000 1158.500000 536.350000 ;
      RECT 382.500000 535.650000 399.000000 536.350000 ;
      RECT 0.000000 535.650000 358.500000 536.350000 ;
      RECT 1166.500000 534.350000 1186.000000 537.650000 ;
      RECT 1157.500000 534.350000 1158.500000 535.650000 ;
      RECT 382.500000 534.350000 383.500000 535.650000 ;
      RECT 366.500000 534.350000 369.500000 537.650000 ;
      RECT 357.500000 534.350000 358.500000 535.650000 ;
      RECT 1157.500000 533.650000 1186.000000 534.350000 ;
      RECT 357.500000 533.650000 383.500000 534.350000 ;
      RECT 1157.500000 532.350000 1158.500000 533.650000 ;
      RECT 1139.000000 532.350000 1149.500000 535.650000 ;
      RECT 396.500000 532.350000 399.000000 535.650000 ;
      RECT 382.500000 532.350000 383.500000 533.650000 ;
      RECT 357.500000 532.350000 358.500000 533.650000 ;
      RECT 0.000000 532.350000 349.500000 535.650000 ;
      RECT 1139.000000 531.650000 1158.500000 532.350000 ;
      RECT 382.500000 531.650000 399.000000 532.350000 ;
      RECT 0.000000 531.650000 358.500000 532.350000 ;
      RECT 1166.500000 530.350000 1186.000000 533.650000 ;
      RECT 1157.500000 530.350000 1158.500000 531.650000 ;
      RECT 382.500000 530.350000 383.500000 531.650000 ;
      RECT 366.500000 530.350000 369.500000 533.650000 ;
      RECT 357.500000 530.350000 358.500000 531.650000 ;
      RECT 1157.500000 529.650000 1186.000000 530.350000 ;
      RECT 357.500000 529.650000 383.500000 530.350000 ;
      RECT 1157.500000 528.350000 1158.500000 529.650000 ;
      RECT 1139.000000 528.350000 1149.500000 531.650000 ;
      RECT 396.500000 528.350000 399.000000 531.650000 ;
      RECT 382.500000 528.350000 383.500000 529.650000 ;
      RECT 357.500000 528.350000 358.500000 529.650000 ;
      RECT 0.000000 528.350000 349.500000 531.650000 ;
      RECT 1139.000000 527.650000 1158.500000 528.350000 ;
      RECT 382.500000 527.650000 399.000000 528.350000 ;
      RECT 0.000000 527.650000 358.500000 528.350000 ;
      RECT 1166.500000 526.350000 1186.000000 529.650000 ;
      RECT 1157.500000 526.350000 1158.500000 527.650000 ;
      RECT 382.500000 526.350000 383.500000 527.650000 ;
      RECT 366.500000 526.350000 369.500000 529.650000 ;
      RECT 357.500000 526.350000 358.500000 527.650000 ;
      RECT 1157.500000 525.650000 1186.000000 526.350000 ;
      RECT 357.500000 525.650000 383.500000 526.350000 ;
      RECT 1157.500000 524.350000 1158.500000 525.650000 ;
      RECT 1139.000000 524.350000 1149.500000 527.650000 ;
      RECT 396.500000 524.350000 399.000000 527.650000 ;
      RECT 382.500000 524.350000 383.500000 525.650000 ;
      RECT 357.500000 524.350000 358.500000 525.650000 ;
      RECT 0.000000 524.350000 349.500000 527.650000 ;
      RECT 1139.000000 523.650000 1158.500000 524.350000 ;
      RECT 382.500000 523.650000 399.000000 524.350000 ;
      RECT 0.000000 523.650000 358.500000 524.350000 ;
      RECT 1166.500000 522.350000 1186.000000 525.650000 ;
      RECT 1157.500000 522.350000 1158.500000 523.650000 ;
      RECT 382.500000 522.350000 383.500000 523.650000 ;
      RECT 366.500000 522.350000 369.500000 525.650000 ;
      RECT 357.500000 522.350000 358.500000 523.650000 ;
      RECT 1157.500000 521.650000 1186.000000 522.350000 ;
      RECT 357.500000 521.650000 383.500000 522.350000 ;
      RECT 1157.500000 520.350000 1158.500000 521.650000 ;
      RECT 1139.000000 520.350000 1149.500000 523.650000 ;
      RECT 396.500000 520.350000 399.000000 523.650000 ;
      RECT 382.500000 520.350000 383.500000 521.650000 ;
      RECT 357.500000 520.350000 358.500000 521.650000 ;
      RECT 0.000000 520.350000 349.500000 523.650000 ;
      RECT 1139.000000 519.650000 1158.500000 520.350000 ;
      RECT 382.500000 519.650000 399.000000 520.350000 ;
      RECT 0.000000 519.650000 358.500000 520.350000 ;
      RECT 1166.500000 518.350000 1186.000000 521.650000 ;
      RECT 1157.500000 518.350000 1158.500000 519.650000 ;
      RECT 382.500000 518.350000 383.500000 519.650000 ;
      RECT 366.500000 518.350000 369.500000 521.650000 ;
      RECT 357.500000 518.350000 358.500000 519.650000 ;
      RECT 1157.500000 517.650000 1186.000000 518.350000 ;
      RECT 357.500000 517.650000 383.500000 518.350000 ;
      RECT 307.500000 517.650000 349.500000 519.650000 ;
      RECT 0.000000 517.650000 299.500000 519.650000 ;
      RECT 1157.500000 516.350000 1158.500000 517.650000 ;
      RECT 1139.000000 516.350000 1149.500000 519.650000 ;
      RECT 396.500000 516.350000 399.000000 519.650000 ;
      RECT 382.500000 516.350000 383.500000 517.650000 ;
      RECT 357.500000 516.350000 358.500000 517.650000 ;
      RECT 316.500000 516.350000 349.500000 517.650000 ;
      RECT 307.500000 516.350000 308.500000 517.650000 ;
      RECT 266.500000 516.350000 299.500000 517.650000 ;
      RECT 1139.000000 515.650000 1158.500000 516.350000 ;
      RECT 382.500000 515.650000 399.000000 516.350000 ;
      RECT 316.500000 515.650000 358.500000 516.350000 ;
      RECT 266.500000 515.650000 308.500000 516.350000 ;
      RECT 216.500000 515.650000 258.500000 517.650000 ;
      RECT 166.500000 515.650000 208.500000 517.650000 ;
      RECT 116.500000 515.650000 158.500000 517.650000 ;
      RECT 66.500000 515.650000 108.500000 517.650000 ;
      RECT 29.500000 515.650000 58.500000 517.650000 ;
      RECT 0.000000 515.650000 16.500000 517.650000 ;
      RECT 1166.500000 514.350000 1186.000000 517.650000 ;
      RECT 1157.500000 514.350000 1158.500000 515.650000 ;
      RECT 382.500000 514.350000 383.500000 515.650000 ;
      RECT 366.500000 514.350000 369.500000 517.650000 ;
      RECT 357.500000 514.350000 358.500000 515.650000 ;
      RECT 316.500000 514.350000 349.500000 515.650000 ;
      RECT 307.500000 514.350000 308.500000 515.650000 ;
      RECT 266.500000 514.350000 299.500000 515.650000 ;
      RECT 257.500000 514.350000 258.500000 515.650000 ;
      RECT 216.500000 514.350000 249.500000 515.650000 ;
      RECT 207.500000 514.350000 208.500000 515.650000 ;
      RECT 166.500000 514.350000 199.500000 515.650000 ;
      RECT 157.500000 514.350000 158.500000 515.650000 ;
      RECT 116.500000 514.350000 149.500000 515.650000 ;
      RECT 107.500000 514.350000 108.500000 515.650000 ;
      RECT 66.500000 514.350000 99.500000 515.650000 ;
      RECT 57.500000 514.350000 58.500000 515.650000 ;
      RECT 29.500000 514.350000 49.500000 515.650000 ;
      RECT 15.500000 514.350000 16.500000 515.650000 ;
      RECT 1157.500000 513.650000 1186.000000 514.350000 ;
      RECT 357.500000 513.650000 383.500000 514.350000 ;
      RECT 307.500000 513.650000 349.500000 514.350000 ;
      RECT 257.500000 513.650000 299.500000 514.350000 ;
      RECT 207.500000 513.650000 249.500000 514.350000 ;
      RECT 157.500000 513.650000 199.500000 514.350000 ;
      RECT 107.500000 513.650000 149.500000 514.350000 ;
      RECT 57.500000 513.650000 99.500000 514.350000 ;
      RECT 15.500000 513.650000 49.500000 514.350000 ;
      RECT 1157.500000 512.350000 1158.500000 513.650000 ;
      RECT 1139.000000 512.350000 1149.500000 515.650000 ;
      RECT 396.500000 512.350000 399.000000 515.650000 ;
      RECT 382.500000 512.350000 383.500000 513.650000 ;
      RECT 357.500000 512.350000 358.500000 513.650000 ;
      RECT 316.500000 512.350000 349.500000 513.650000 ;
      RECT 307.500000 512.350000 308.500000 513.650000 ;
      RECT 266.500000 512.350000 299.500000 513.650000 ;
      RECT 257.500000 512.350000 258.500000 513.650000 ;
      RECT 216.500000 512.350000 249.500000 513.650000 ;
      RECT 207.500000 512.350000 208.500000 513.650000 ;
      RECT 166.500000 512.350000 199.500000 513.650000 ;
      RECT 157.500000 512.350000 158.500000 513.650000 ;
      RECT 116.500000 512.350000 149.500000 513.650000 ;
      RECT 107.500000 512.350000 108.500000 513.650000 ;
      RECT 66.500000 512.350000 99.500000 513.650000 ;
      RECT 57.500000 512.350000 58.500000 513.650000 ;
      RECT 29.500000 512.350000 49.500000 513.650000 ;
      RECT 15.500000 512.350000 16.500000 513.650000 ;
      RECT 0.000000 512.350000 2.500000 515.650000 ;
      RECT 1139.000000 511.650000 1158.500000 512.350000 ;
      RECT 382.500000 511.650000 399.000000 512.350000 ;
      RECT 316.500000 511.650000 358.500000 512.350000 ;
      RECT 266.500000 511.650000 308.500000 512.350000 ;
      RECT 216.500000 511.650000 258.500000 512.350000 ;
      RECT 166.500000 511.650000 208.500000 512.350000 ;
      RECT 116.500000 511.650000 158.500000 512.350000 ;
      RECT 66.500000 511.650000 108.500000 512.350000 ;
      RECT 29.500000 511.650000 58.500000 512.350000 ;
      RECT 0.000000 511.650000 16.500000 512.350000 ;
      RECT 1166.500000 510.350000 1186.000000 513.650000 ;
      RECT 1157.500000 510.350000 1158.500000 511.650000 ;
      RECT 382.500000 510.350000 383.500000 511.650000 ;
      RECT 366.500000 510.350000 369.500000 513.650000 ;
      RECT 357.500000 510.350000 358.500000 511.650000 ;
      RECT 316.500000 510.350000 349.500000 511.650000 ;
      RECT 307.500000 510.350000 308.500000 511.650000 ;
      RECT 266.500000 510.350000 299.500000 511.650000 ;
      RECT 257.500000 510.350000 258.500000 511.650000 ;
      RECT 216.500000 510.350000 249.500000 511.650000 ;
      RECT 207.500000 510.350000 208.500000 511.650000 ;
      RECT 166.500000 510.350000 199.500000 511.650000 ;
      RECT 157.500000 510.350000 158.500000 511.650000 ;
      RECT 116.500000 510.350000 149.500000 511.650000 ;
      RECT 107.500000 510.350000 108.500000 511.650000 ;
      RECT 66.500000 510.350000 99.500000 511.650000 ;
      RECT 57.500000 510.350000 58.500000 511.650000 ;
      RECT 29.500000 510.350000 49.500000 511.650000 ;
      RECT 15.500000 510.350000 16.500000 511.650000 ;
      RECT 1157.500000 509.650000 1186.000000 510.350000 ;
      RECT 357.500000 509.650000 383.500000 510.350000 ;
      RECT 307.500000 509.650000 349.500000 510.350000 ;
      RECT 257.500000 509.650000 299.500000 510.350000 ;
      RECT 207.500000 509.650000 249.500000 510.350000 ;
      RECT 157.500000 509.650000 199.500000 510.350000 ;
      RECT 107.500000 509.650000 149.500000 510.350000 ;
      RECT 57.500000 509.650000 99.500000 510.350000 ;
      RECT 15.500000 509.650000 49.500000 510.350000 ;
      RECT 1157.500000 508.350000 1158.500000 509.650000 ;
      RECT 1139.000000 508.350000 1149.500000 511.650000 ;
      RECT 396.500000 508.350000 399.000000 511.650000 ;
      RECT 382.500000 508.350000 383.500000 509.650000 ;
      RECT 357.500000 508.350000 358.500000 509.650000 ;
      RECT 316.500000 508.350000 349.500000 509.650000 ;
      RECT 307.500000 508.350000 308.500000 509.650000 ;
      RECT 266.500000 508.350000 299.500000 509.650000 ;
      RECT 257.500000 508.350000 258.500000 509.650000 ;
      RECT 216.500000 508.350000 249.500000 509.650000 ;
      RECT 207.500000 508.350000 208.500000 509.650000 ;
      RECT 166.500000 508.350000 199.500000 509.650000 ;
      RECT 157.500000 508.350000 158.500000 509.650000 ;
      RECT 116.500000 508.350000 149.500000 509.650000 ;
      RECT 107.500000 508.350000 108.500000 509.650000 ;
      RECT 66.500000 508.350000 99.500000 509.650000 ;
      RECT 57.500000 508.350000 58.500000 509.650000 ;
      RECT 29.500000 508.350000 49.500000 509.650000 ;
      RECT 15.500000 508.350000 16.500000 509.650000 ;
      RECT 0.000000 508.350000 2.500000 511.650000 ;
      RECT 1139.000000 507.650000 1158.500000 508.350000 ;
      RECT 382.500000 507.650000 399.000000 508.350000 ;
      RECT 316.500000 507.650000 358.500000 508.350000 ;
      RECT 266.500000 507.650000 308.500000 508.350000 ;
      RECT 216.500000 507.650000 258.500000 508.350000 ;
      RECT 166.500000 507.650000 208.500000 508.350000 ;
      RECT 116.500000 507.650000 158.500000 508.350000 ;
      RECT 66.500000 507.650000 108.500000 508.350000 ;
      RECT 29.500000 507.650000 58.500000 508.350000 ;
      RECT 0.000000 507.650000 16.500000 508.350000 ;
      RECT 1166.500000 506.350000 1186.000000 509.650000 ;
      RECT 1157.500000 506.350000 1158.500000 507.650000 ;
      RECT 382.500000 506.350000 383.500000 507.650000 ;
      RECT 366.500000 506.350000 369.500000 509.650000 ;
      RECT 357.500000 506.350000 358.500000 507.650000 ;
      RECT 316.500000 506.350000 349.500000 507.650000 ;
      RECT 307.500000 506.350000 308.500000 507.650000 ;
      RECT 266.500000 506.350000 299.500000 507.650000 ;
      RECT 257.500000 506.350000 258.500000 507.650000 ;
      RECT 216.500000 506.350000 249.500000 507.650000 ;
      RECT 207.500000 506.350000 208.500000 507.650000 ;
      RECT 166.500000 506.350000 199.500000 507.650000 ;
      RECT 157.500000 506.350000 158.500000 507.650000 ;
      RECT 116.500000 506.350000 149.500000 507.650000 ;
      RECT 107.500000 506.350000 108.500000 507.650000 ;
      RECT 66.500000 506.350000 99.500000 507.650000 ;
      RECT 57.500000 506.350000 58.500000 507.650000 ;
      RECT 29.500000 506.350000 49.500000 507.650000 ;
      RECT 15.500000 506.350000 16.500000 507.650000 ;
      RECT 396.500000 506.000000 399.000000 507.650000 ;
      RECT 1157.500000 505.650000 1186.000000 506.350000 ;
      RECT 396.500000 505.650000 749.000000 506.000000 ;
      RECT 357.500000 505.650000 383.500000 506.350000 ;
      RECT 307.500000 505.650000 349.500000 506.350000 ;
      RECT 257.500000 505.650000 299.500000 506.350000 ;
      RECT 207.500000 505.650000 249.500000 506.350000 ;
      RECT 157.500000 505.650000 199.500000 506.350000 ;
      RECT 107.500000 505.650000 149.500000 506.350000 ;
      RECT 57.500000 505.650000 99.500000 506.350000 ;
      RECT 15.500000 505.650000 49.500000 506.350000 ;
      RECT 1157.500000 504.350000 1158.500000 505.650000 ;
      RECT 1139.000000 504.350000 1149.500000 507.650000 ;
      RECT 396.500000 504.350000 408.500000 505.650000 ;
      RECT 382.500000 504.350000 383.500000 505.650000 ;
      RECT 357.500000 504.350000 358.500000 505.650000 ;
      RECT 316.500000 504.350000 349.500000 505.650000 ;
      RECT 307.500000 504.350000 308.500000 505.650000 ;
      RECT 266.500000 504.350000 299.500000 505.650000 ;
      RECT 257.500000 504.350000 258.500000 505.650000 ;
      RECT 216.500000 504.350000 249.500000 505.650000 ;
      RECT 207.500000 504.350000 208.500000 505.650000 ;
      RECT 166.500000 504.350000 199.500000 505.650000 ;
      RECT 157.500000 504.350000 158.500000 505.650000 ;
      RECT 116.500000 504.350000 149.500000 505.650000 ;
      RECT 107.500000 504.350000 108.500000 505.650000 ;
      RECT 66.500000 504.350000 99.500000 505.650000 ;
      RECT 57.500000 504.350000 58.500000 505.650000 ;
      RECT 29.500000 504.350000 49.500000 505.650000 ;
      RECT 15.500000 504.350000 16.500000 505.650000 ;
      RECT 0.000000 504.350000 2.500000 507.650000 ;
      RECT 1139.000000 503.650000 1158.500000 504.350000 ;
      RECT 716.500000 503.650000 749.000000 505.650000 ;
      RECT 666.500000 503.650000 708.500000 505.650000 ;
      RECT 616.500000 503.650000 658.500000 505.650000 ;
      RECT 566.500000 503.650000 608.500000 505.650000 ;
      RECT 516.500000 503.650000 558.500000 505.650000 ;
      RECT 466.500000 503.650000 508.500000 505.650000 ;
      RECT 416.500000 503.650000 458.500000 505.650000 ;
      RECT 382.500000 503.650000 408.500000 504.350000 ;
      RECT 316.500000 503.650000 358.500000 504.350000 ;
      RECT 266.500000 503.650000 308.500000 504.350000 ;
      RECT 216.500000 503.650000 258.500000 504.350000 ;
      RECT 166.500000 503.650000 208.500000 504.350000 ;
      RECT 116.500000 503.650000 158.500000 504.350000 ;
      RECT 66.500000 503.650000 108.500000 504.350000 ;
      RECT 29.500000 503.650000 58.500000 504.350000 ;
      RECT 0.000000 503.650000 16.500000 504.350000 ;
      RECT 1166.500000 502.350000 1186.000000 505.650000 ;
      RECT 1157.500000 502.350000 1158.500000 503.650000 ;
      RECT 716.500000 502.350000 733.500000 503.650000 ;
      RECT 707.500000 502.350000 708.500000 503.650000 ;
      RECT 666.500000 502.350000 699.500000 503.650000 ;
      RECT 657.500000 502.350000 658.500000 503.650000 ;
      RECT 616.500000 502.350000 649.500000 503.650000 ;
      RECT 607.500000 502.350000 608.500000 503.650000 ;
      RECT 566.500000 502.350000 599.500000 503.650000 ;
      RECT 557.500000 502.350000 558.500000 503.650000 ;
      RECT 516.500000 502.350000 549.500000 503.650000 ;
      RECT 507.500000 502.350000 508.500000 503.650000 ;
      RECT 466.500000 502.350000 499.500000 503.650000 ;
      RECT 457.500000 502.350000 458.500000 503.650000 ;
      RECT 416.500000 502.350000 449.500000 503.650000 ;
      RECT 407.500000 502.350000 408.500000 503.650000 ;
      RECT 382.500000 502.350000 383.500000 503.650000 ;
      RECT 366.500000 502.350000 369.500000 505.650000 ;
      RECT 357.500000 502.350000 358.500000 503.650000 ;
      RECT 316.500000 502.350000 349.500000 503.650000 ;
      RECT 307.500000 502.350000 308.500000 503.650000 ;
      RECT 266.500000 502.350000 299.500000 503.650000 ;
      RECT 257.500000 502.350000 258.500000 503.650000 ;
      RECT 216.500000 502.350000 249.500000 503.650000 ;
      RECT 207.500000 502.350000 208.500000 503.650000 ;
      RECT 166.500000 502.350000 199.500000 503.650000 ;
      RECT 157.500000 502.350000 158.500000 503.650000 ;
      RECT 116.500000 502.350000 149.500000 503.650000 ;
      RECT 107.500000 502.350000 108.500000 503.650000 ;
      RECT 66.500000 502.350000 99.500000 503.650000 ;
      RECT 57.500000 502.350000 58.500000 503.650000 ;
      RECT 29.500000 502.350000 49.500000 503.650000 ;
      RECT 15.500000 502.350000 16.500000 503.650000 ;
      RECT 1157.500000 501.650000 1186.000000 502.350000 ;
      RECT 707.500000 501.650000 733.500000 502.350000 ;
      RECT 657.500000 501.650000 699.500000 502.350000 ;
      RECT 607.500000 501.650000 649.500000 502.350000 ;
      RECT 557.500000 501.650000 599.500000 502.350000 ;
      RECT 507.500000 501.650000 549.500000 502.350000 ;
      RECT 457.500000 501.650000 499.500000 502.350000 ;
      RECT 407.500000 501.650000 449.500000 502.350000 ;
      RECT 357.500000 501.650000 383.500000 502.350000 ;
      RECT 307.500000 501.650000 349.500000 502.350000 ;
      RECT 257.500000 501.650000 299.500000 502.350000 ;
      RECT 207.500000 501.650000 249.500000 502.350000 ;
      RECT 157.500000 501.650000 199.500000 502.350000 ;
      RECT 107.500000 501.650000 149.500000 502.350000 ;
      RECT 57.500000 501.650000 99.500000 502.350000 ;
      RECT 15.500000 501.650000 49.500000 502.350000 ;
      RECT 1157.500000 500.350000 1158.500000 501.650000 ;
      RECT 1139.000000 500.350000 1149.500000 503.650000 ;
      RECT 746.500000 500.350000 749.000000 503.650000 ;
      RECT 716.500000 500.350000 733.500000 501.650000 ;
      RECT 707.500000 500.350000 708.500000 501.650000 ;
      RECT 666.500000 500.350000 699.500000 501.650000 ;
      RECT 657.500000 500.350000 658.500000 501.650000 ;
      RECT 616.500000 500.350000 649.500000 501.650000 ;
      RECT 607.500000 500.350000 608.500000 501.650000 ;
      RECT 566.500000 500.350000 599.500000 501.650000 ;
      RECT 557.500000 500.350000 558.500000 501.650000 ;
      RECT 516.500000 500.350000 549.500000 501.650000 ;
      RECT 507.500000 500.350000 508.500000 501.650000 ;
      RECT 466.500000 500.350000 499.500000 501.650000 ;
      RECT 457.500000 500.350000 458.500000 501.650000 ;
      RECT 416.500000 500.350000 449.500000 501.650000 ;
      RECT 407.500000 500.350000 408.500000 501.650000 ;
      RECT 396.500000 500.350000 399.500000 503.650000 ;
      RECT 382.500000 500.350000 383.500000 501.650000 ;
      RECT 357.500000 500.350000 358.500000 501.650000 ;
      RECT 316.500000 500.350000 349.500000 501.650000 ;
      RECT 307.500000 500.350000 308.500000 501.650000 ;
      RECT 266.500000 500.350000 299.500000 501.650000 ;
      RECT 257.500000 500.350000 258.500000 501.650000 ;
      RECT 216.500000 500.350000 249.500000 501.650000 ;
      RECT 207.500000 500.350000 208.500000 501.650000 ;
      RECT 166.500000 500.350000 199.500000 501.650000 ;
      RECT 157.500000 500.350000 158.500000 501.650000 ;
      RECT 116.500000 500.350000 149.500000 501.650000 ;
      RECT 107.500000 500.350000 108.500000 501.650000 ;
      RECT 66.500000 500.350000 99.500000 501.650000 ;
      RECT 57.500000 500.350000 58.500000 501.650000 ;
      RECT 29.500000 500.350000 49.500000 501.650000 ;
      RECT 15.500000 500.350000 16.500000 501.650000 ;
      RECT 0.000000 500.350000 2.500000 503.650000 ;
      RECT 1139.000000 499.650000 1158.500000 500.350000 ;
      RECT 716.500000 499.650000 749.000000 500.350000 ;
      RECT 666.500000 499.650000 708.500000 500.350000 ;
      RECT 616.500000 499.650000 658.500000 500.350000 ;
      RECT 566.500000 499.650000 608.500000 500.350000 ;
      RECT 516.500000 499.650000 558.500000 500.350000 ;
      RECT 466.500000 499.650000 508.500000 500.350000 ;
      RECT 416.500000 499.650000 458.500000 500.350000 ;
      RECT 382.500000 499.650000 408.500000 500.350000 ;
      RECT 316.500000 499.650000 358.500000 500.350000 ;
      RECT 266.500000 499.650000 308.500000 500.350000 ;
      RECT 216.500000 499.650000 258.500000 500.350000 ;
      RECT 166.500000 499.650000 208.500000 500.350000 ;
      RECT 116.500000 499.650000 158.500000 500.350000 ;
      RECT 66.500000 499.650000 108.500000 500.350000 ;
      RECT 29.500000 499.650000 58.500000 500.350000 ;
      RECT 0.000000 499.650000 16.500000 500.350000 ;
      RECT 1166.500000 498.350000 1186.000000 501.650000 ;
      RECT 1157.500000 498.350000 1158.500000 499.650000 ;
      RECT 716.500000 498.350000 733.500000 499.650000 ;
      RECT 707.500000 498.350000 708.500000 499.650000 ;
      RECT 666.500000 498.350000 699.500000 499.650000 ;
      RECT 657.500000 498.350000 658.500000 499.650000 ;
      RECT 616.500000 498.350000 649.500000 499.650000 ;
      RECT 607.500000 498.350000 608.500000 499.650000 ;
      RECT 566.500000 498.350000 599.500000 499.650000 ;
      RECT 557.500000 498.350000 558.500000 499.650000 ;
      RECT 516.500000 498.350000 549.500000 499.650000 ;
      RECT 507.500000 498.350000 508.500000 499.650000 ;
      RECT 466.500000 498.350000 499.500000 499.650000 ;
      RECT 457.500000 498.350000 458.500000 499.650000 ;
      RECT 416.500000 498.350000 449.500000 499.650000 ;
      RECT 407.500000 498.350000 408.500000 499.650000 ;
      RECT 382.500000 498.350000 383.500000 499.650000 ;
      RECT 366.500000 498.350000 369.500000 501.650000 ;
      RECT 357.500000 498.350000 358.500000 499.650000 ;
      RECT 316.500000 498.350000 349.500000 499.650000 ;
      RECT 307.500000 498.350000 308.500000 499.650000 ;
      RECT 266.500000 498.350000 299.500000 499.650000 ;
      RECT 257.500000 498.350000 258.500000 499.650000 ;
      RECT 216.500000 498.350000 249.500000 499.650000 ;
      RECT 207.500000 498.350000 208.500000 499.650000 ;
      RECT 166.500000 498.350000 199.500000 499.650000 ;
      RECT 157.500000 498.350000 158.500000 499.650000 ;
      RECT 116.500000 498.350000 149.500000 499.650000 ;
      RECT 107.500000 498.350000 108.500000 499.650000 ;
      RECT 66.500000 498.350000 99.500000 499.650000 ;
      RECT 57.500000 498.350000 58.500000 499.650000 ;
      RECT 29.500000 498.350000 49.500000 499.650000 ;
      RECT 15.500000 498.350000 16.500000 499.650000 ;
      RECT 1157.500000 497.650000 1186.000000 498.350000 ;
      RECT 707.500000 497.650000 733.500000 498.350000 ;
      RECT 657.500000 497.650000 699.500000 498.350000 ;
      RECT 607.500000 497.650000 649.500000 498.350000 ;
      RECT 557.500000 497.650000 599.500000 498.350000 ;
      RECT 507.500000 497.650000 549.500000 498.350000 ;
      RECT 457.500000 497.650000 499.500000 498.350000 ;
      RECT 407.500000 497.650000 449.500000 498.350000 ;
      RECT 357.500000 497.650000 383.500000 498.350000 ;
      RECT 307.500000 497.650000 349.500000 498.350000 ;
      RECT 257.500000 497.650000 299.500000 498.350000 ;
      RECT 207.500000 497.650000 249.500000 498.350000 ;
      RECT 157.500000 497.650000 199.500000 498.350000 ;
      RECT 107.500000 497.650000 149.500000 498.350000 ;
      RECT 57.500000 497.650000 99.500000 498.350000 ;
      RECT 15.500000 497.650000 49.500000 498.350000 ;
      RECT 1157.500000 496.350000 1158.500000 497.650000 ;
      RECT 1139.000000 496.350000 1149.500000 499.650000 ;
      RECT 746.500000 496.350000 749.000000 499.650000 ;
      RECT 716.500000 496.350000 733.500000 497.650000 ;
      RECT 707.500000 496.350000 708.500000 497.650000 ;
      RECT 666.500000 496.350000 699.500000 497.650000 ;
      RECT 657.500000 496.350000 658.500000 497.650000 ;
      RECT 616.500000 496.350000 649.500000 497.650000 ;
      RECT 607.500000 496.350000 608.500000 497.650000 ;
      RECT 566.500000 496.350000 599.500000 497.650000 ;
      RECT 557.500000 496.350000 558.500000 497.650000 ;
      RECT 516.500000 496.350000 549.500000 497.650000 ;
      RECT 507.500000 496.350000 508.500000 497.650000 ;
      RECT 466.500000 496.350000 499.500000 497.650000 ;
      RECT 457.500000 496.350000 458.500000 497.650000 ;
      RECT 416.500000 496.350000 449.500000 497.650000 ;
      RECT 407.500000 496.350000 408.500000 497.650000 ;
      RECT 396.500000 496.350000 399.500000 499.650000 ;
      RECT 382.500000 496.350000 383.500000 497.650000 ;
      RECT 357.500000 496.350000 358.500000 497.650000 ;
      RECT 316.500000 496.350000 349.500000 497.650000 ;
      RECT 307.500000 496.350000 308.500000 497.650000 ;
      RECT 266.500000 496.350000 299.500000 497.650000 ;
      RECT 257.500000 496.350000 258.500000 497.650000 ;
      RECT 216.500000 496.350000 249.500000 497.650000 ;
      RECT 207.500000 496.350000 208.500000 497.650000 ;
      RECT 166.500000 496.350000 199.500000 497.650000 ;
      RECT 157.500000 496.350000 158.500000 497.650000 ;
      RECT 116.500000 496.350000 149.500000 497.650000 ;
      RECT 107.500000 496.350000 108.500000 497.650000 ;
      RECT 66.500000 496.350000 99.500000 497.650000 ;
      RECT 57.500000 496.350000 58.500000 497.650000 ;
      RECT 29.500000 496.350000 49.500000 497.650000 ;
      RECT 15.500000 496.350000 16.500000 497.650000 ;
      RECT 0.000000 496.350000 2.500000 499.650000 ;
      RECT 1139.000000 495.650000 1158.500000 496.350000 ;
      RECT 716.500000 495.650000 749.000000 496.350000 ;
      RECT 666.500000 495.650000 708.500000 496.350000 ;
      RECT 616.500000 495.650000 658.500000 496.350000 ;
      RECT 566.500000 495.650000 608.500000 496.350000 ;
      RECT 516.500000 495.650000 558.500000 496.350000 ;
      RECT 466.500000 495.650000 508.500000 496.350000 ;
      RECT 416.500000 495.650000 458.500000 496.350000 ;
      RECT 382.500000 495.650000 408.500000 496.350000 ;
      RECT 316.500000 495.650000 358.500000 496.350000 ;
      RECT 266.500000 495.650000 308.500000 496.350000 ;
      RECT 216.500000 495.650000 258.500000 496.350000 ;
      RECT 166.500000 495.650000 208.500000 496.350000 ;
      RECT 116.500000 495.650000 158.500000 496.350000 ;
      RECT 66.500000 495.650000 108.500000 496.350000 ;
      RECT 29.500000 495.650000 58.500000 496.350000 ;
      RECT 0.000000 495.650000 16.500000 496.350000 ;
      RECT 1166.500000 494.350000 1186.000000 497.650000 ;
      RECT 1157.500000 494.350000 1158.500000 495.650000 ;
      RECT 716.500000 494.350000 733.500000 495.650000 ;
      RECT 707.500000 494.350000 708.500000 495.650000 ;
      RECT 666.500000 494.350000 699.500000 495.650000 ;
      RECT 657.500000 494.350000 658.500000 495.650000 ;
      RECT 616.500000 494.350000 649.500000 495.650000 ;
      RECT 607.500000 494.350000 608.500000 495.650000 ;
      RECT 566.500000 494.350000 599.500000 495.650000 ;
      RECT 557.500000 494.350000 558.500000 495.650000 ;
      RECT 516.500000 494.350000 549.500000 495.650000 ;
      RECT 507.500000 494.350000 508.500000 495.650000 ;
      RECT 466.500000 494.350000 499.500000 495.650000 ;
      RECT 457.500000 494.350000 458.500000 495.650000 ;
      RECT 416.500000 494.350000 449.500000 495.650000 ;
      RECT 407.500000 494.350000 408.500000 495.650000 ;
      RECT 382.500000 494.350000 383.500000 495.650000 ;
      RECT 366.500000 494.350000 369.500000 497.650000 ;
      RECT 357.500000 494.350000 358.500000 495.650000 ;
      RECT 316.500000 494.350000 349.500000 495.650000 ;
      RECT 307.500000 494.350000 308.500000 495.650000 ;
      RECT 266.500000 494.350000 299.500000 495.650000 ;
      RECT 257.500000 494.350000 258.500000 495.650000 ;
      RECT 216.500000 494.350000 249.500000 495.650000 ;
      RECT 207.500000 494.350000 208.500000 495.650000 ;
      RECT 166.500000 494.350000 199.500000 495.650000 ;
      RECT 157.500000 494.350000 158.500000 495.650000 ;
      RECT 116.500000 494.350000 149.500000 495.650000 ;
      RECT 107.500000 494.350000 108.500000 495.650000 ;
      RECT 66.500000 494.350000 99.500000 495.650000 ;
      RECT 57.500000 494.350000 58.500000 495.650000 ;
      RECT 29.500000 494.350000 49.500000 495.650000 ;
      RECT 15.500000 494.350000 16.500000 495.650000 ;
      RECT 1157.500000 493.650000 1186.000000 494.350000 ;
      RECT 707.500000 493.650000 733.500000 494.350000 ;
      RECT 657.500000 493.650000 699.500000 494.350000 ;
      RECT 607.500000 493.650000 649.500000 494.350000 ;
      RECT 557.500000 493.650000 599.500000 494.350000 ;
      RECT 507.500000 493.650000 549.500000 494.350000 ;
      RECT 457.500000 493.650000 499.500000 494.350000 ;
      RECT 407.500000 493.650000 449.500000 494.350000 ;
      RECT 357.500000 493.650000 383.500000 494.350000 ;
      RECT 307.500000 493.650000 349.500000 494.350000 ;
      RECT 257.500000 493.650000 299.500000 494.350000 ;
      RECT 207.500000 493.650000 249.500000 494.350000 ;
      RECT 157.500000 493.650000 199.500000 494.350000 ;
      RECT 107.500000 493.650000 149.500000 494.350000 ;
      RECT 57.500000 493.650000 99.500000 494.350000 ;
      RECT 15.500000 493.650000 49.500000 494.350000 ;
      RECT 1157.500000 492.350000 1158.500000 493.650000 ;
      RECT 1139.000000 492.350000 1149.500000 495.650000 ;
      RECT 746.500000 492.350000 749.000000 495.650000 ;
      RECT 716.500000 492.350000 733.500000 493.650000 ;
      RECT 707.500000 492.350000 708.500000 493.650000 ;
      RECT 666.500000 492.350000 699.500000 493.650000 ;
      RECT 657.500000 492.350000 658.500000 493.650000 ;
      RECT 616.500000 492.350000 649.500000 493.650000 ;
      RECT 607.500000 492.350000 608.500000 493.650000 ;
      RECT 566.500000 492.350000 599.500000 493.650000 ;
      RECT 557.500000 492.350000 558.500000 493.650000 ;
      RECT 516.500000 492.350000 549.500000 493.650000 ;
      RECT 507.500000 492.350000 508.500000 493.650000 ;
      RECT 466.500000 492.350000 499.500000 493.650000 ;
      RECT 457.500000 492.350000 458.500000 493.650000 ;
      RECT 416.500000 492.350000 449.500000 493.650000 ;
      RECT 407.500000 492.350000 408.500000 493.650000 ;
      RECT 396.500000 492.350000 399.500000 495.650000 ;
      RECT 382.500000 492.350000 383.500000 493.650000 ;
      RECT 357.500000 492.350000 358.500000 493.650000 ;
      RECT 316.500000 492.350000 349.500000 493.650000 ;
      RECT 307.500000 492.350000 308.500000 493.650000 ;
      RECT 266.500000 492.350000 299.500000 493.650000 ;
      RECT 257.500000 492.350000 258.500000 493.650000 ;
      RECT 216.500000 492.350000 249.500000 493.650000 ;
      RECT 207.500000 492.350000 208.500000 493.650000 ;
      RECT 166.500000 492.350000 199.500000 493.650000 ;
      RECT 157.500000 492.350000 158.500000 493.650000 ;
      RECT 116.500000 492.350000 149.500000 493.650000 ;
      RECT 107.500000 492.350000 108.500000 493.650000 ;
      RECT 66.500000 492.350000 99.500000 493.650000 ;
      RECT 57.500000 492.350000 58.500000 493.650000 ;
      RECT 29.500000 492.350000 49.500000 493.650000 ;
      RECT 15.500000 492.350000 16.500000 493.650000 ;
      RECT 0.000000 492.350000 2.500000 495.650000 ;
      RECT 1139.000000 491.650000 1158.500000 492.350000 ;
      RECT 716.500000 491.650000 749.000000 492.350000 ;
      RECT 666.500000 491.650000 708.500000 492.350000 ;
      RECT 616.500000 491.650000 658.500000 492.350000 ;
      RECT 566.500000 491.650000 608.500000 492.350000 ;
      RECT 516.500000 491.650000 558.500000 492.350000 ;
      RECT 466.500000 491.650000 508.500000 492.350000 ;
      RECT 416.500000 491.650000 458.500000 492.350000 ;
      RECT 382.500000 491.650000 408.500000 492.350000 ;
      RECT 316.500000 491.650000 358.500000 492.350000 ;
      RECT 266.500000 491.650000 308.500000 492.350000 ;
      RECT 216.500000 491.650000 258.500000 492.350000 ;
      RECT 166.500000 491.650000 208.500000 492.350000 ;
      RECT 116.500000 491.650000 158.500000 492.350000 ;
      RECT 66.500000 491.650000 108.500000 492.350000 ;
      RECT 29.500000 491.650000 58.500000 492.350000 ;
      RECT 0.000000 491.650000 16.500000 492.350000 ;
      RECT 1166.500000 490.350000 1186.000000 493.650000 ;
      RECT 1157.500000 490.350000 1158.500000 491.650000 ;
      RECT 716.500000 490.350000 733.500000 491.650000 ;
      RECT 707.500000 490.350000 708.500000 491.650000 ;
      RECT 666.500000 490.350000 699.500000 491.650000 ;
      RECT 657.500000 490.350000 658.500000 491.650000 ;
      RECT 616.500000 490.350000 649.500000 491.650000 ;
      RECT 607.500000 490.350000 608.500000 491.650000 ;
      RECT 566.500000 490.350000 599.500000 491.650000 ;
      RECT 557.500000 490.350000 558.500000 491.650000 ;
      RECT 516.500000 490.350000 549.500000 491.650000 ;
      RECT 507.500000 490.350000 508.500000 491.650000 ;
      RECT 466.500000 490.350000 499.500000 491.650000 ;
      RECT 457.500000 490.350000 458.500000 491.650000 ;
      RECT 416.500000 490.350000 449.500000 491.650000 ;
      RECT 407.500000 490.350000 408.500000 491.650000 ;
      RECT 382.500000 490.350000 399.500000 491.650000 ;
      RECT 366.500000 490.350000 369.500000 493.650000 ;
      RECT 357.500000 490.350000 358.500000 491.650000 ;
      RECT 316.500000 490.350000 349.500000 491.650000 ;
      RECT 307.500000 490.350000 308.500000 491.650000 ;
      RECT 266.500000 490.350000 299.500000 491.650000 ;
      RECT 257.500000 490.350000 258.500000 491.650000 ;
      RECT 216.500000 490.350000 249.500000 491.650000 ;
      RECT 207.500000 490.350000 208.500000 491.650000 ;
      RECT 166.500000 490.350000 199.500000 491.650000 ;
      RECT 157.500000 490.350000 158.500000 491.650000 ;
      RECT 116.500000 490.350000 149.500000 491.650000 ;
      RECT 107.500000 490.350000 108.500000 491.650000 ;
      RECT 66.500000 490.350000 99.500000 491.650000 ;
      RECT 57.500000 490.350000 58.500000 491.650000 ;
      RECT 29.500000 490.350000 49.500000 491.650000 ;
      RECT 15.500000 490.350000 16.500000 491.650000 ;
      RECT 1157.500000 489.650000 1186.000000 490.350000 ;
      RECT 707.500000 489.650000 733.500000 490.350000 ;
      RECT 657.500000 489.650000 699.500000 490.350000 ;
      RECT 607.500000 489.650000 649.500000 490.350000 ;
      RECT 557.500000 489.650000 599.500000 490.350000 ;
      RECT 507.500000 489.650000 549.500000 490.350000 ;
      RECT 457.500000 489.650000 499.500000 490.350000 ;
      RECT 407.500000 489.650000 449.500000 490.350000 ;
      RECT 357.500000 489.650000 399.500000 490.350000 ;
      RECT 307.500000 489.650000 349.500000 490.350000 ;
      RECT 257.500000 489.650000 299.500000 490.350000 ;
      RECT 207.500000 489.650000 249.500000 490.350000 ;
      RECT 157.500000 489.650000 199.500000 490.350000 ;
      RECT 107.500000 489.650000 149.500000 490.350000 ;
      RECT 57.500000 489.650000 99.500000 490.350000 ;
      RECT 15.500000 489.650000 49.500000 490.350000 ;
      RECT 1157.500000 488.350000 1158.500000 489.650000 ;
      RECT 1139.000000 488.350000 1149.500000 491.650000 ;
      RECT 746.500000 488.350000 749.000000 491.650000 ;
      RECT 732.500000 488.350000 733.500000 489.650000 ;
      RECT 707.500000 488.350000 708.500000 489.650000 ;
      RECT 666.500000 488.350000 699.500000 489.650000 ;
      RECT 657.500000 488.350000 658.500000 489.650000 ;
      RECT 616.500000 488.350000 649.500000 489.650000 ;
      RECT 607.500000 488.350000 608.500000 489.650000 ;
      RECT 566.500000 488.350000 599.500000 489.650000 ;
      RECT 557.500000 488.350000 558.500000 489.650000 ;
      RECT 516.500000 488.350000 549.500000 489.650000 ;
      RECT 507.500000 488.350000 508.500000 489.650000 ;
      RECT 466.500000 488.350000 499.500000 489.650000 ;
      RECT 457.500000 488.350000 458.500000 489.650000 ;
      RECT 416.500000 488.350000 449.500000 489.650000 ;
      RECT 407.500000 488.350000 408.500000 489.650000 ;
      RECT 382.500000 488.350000 399.500000 489.650000 ;
      RECT 357.500000 488.350000 358.500000 489.650000 ;
      RECT 316.500000 488.350000 349.500000 489.650000 ;
      RECT 307.500000 488.350000 308.500000 489.650000 ;
      RECT 266.500000 488.350000 299.500000 489.650000 ;
      RECT 257.500000 488.350000 258.500000 489.650000 ;
      RECT 216.500000 488.350000 249.500000 489.650000 ;
      RECT 207.500000 488.350000 208.500000 489.650000 ;
      RECT 166.500000 488.350000 199.500000 489.650000 ;
      RECT 157.500000 488.350000 158.500000 489.650000 ;
      RECT 116.500000 488.350000 149.500000 489.650000 ;
      RECT 107.500000 488.350000 108.500000 489.650000 ;
      RECT 66.500000 488.350000 99.500000 489.650000 ;
      RECT 57.500000 488.350000 58.500000 489.650000 ;
      RECT 29.500000 488.350000 49.500000 489.650000 ;
      RECT 15.500000 488.350000 16.500000 489.650000 ;
      RECT 0.000000 488.350000 2.500000 491.650000 ;
      RECT 1139.000000 487.650000 1158.500000 488.350000 ;
      RECT 732.500000 487.650000 749.000000 488.350000 ;
      RECT 666.500000 487.650000 708.500000 488.350000 ;
      RECT 616.500000 487.650000 658.500000 488.350000 ;
      RECT 566.500000 487.650000 608.500000 488.350000 ;
      RECT 516.500000 487.650000 558.500000 488.350000 ;
      RECT 466.500000 487.650000 508.500000 488.350000 ;
      RECT 416.500000 487.650000 458.500000 488.350000 ;
      RECT 382.500000 487.650000 408.500000 488.350000 ;
      RECT 316.500000 487.650000 358.500000 488.350000 ;
      RECT 266.500000 487.650000 308.500000 488.350000 ;
      RECT 216.500000 487.650000 258.500000 488.350000 ;
      RECT 166.500000 487.650000 208.500000 488.350000 ;
      RECT 116.500000 487.650000 158.500000 488.350000 ;
      RECT 66.500000 487.650000 108.500000 488.350000 ;
      RECT 29.500000 487.650000 58.500000 488.350000 ;
      RECT 0.000000 487.650000 16.500000 488.350000 ;
      RECT 0.000000 487.170000 2.500000 487.650000 ;
      RECT 1166.500000 487.165000 1186.000000 489.650000 ;
      RECT 1166.500000 486.350000 1183.980000 487.165000 ;
      RECT 1157.500000 486.350000 1158.500000 487.650000 ;
      RECT 732.500000 486.350000 733.500000 487.650000 ;
      RECT 716.500000 486.350000 719.500000 489.650000 ;
      RECT 707.500000 486.350000 708.500000 487.650000 ;
      RECT 666.500000 486.350000 699.500000 487.650000 ;
      RECT 657.500000 486.350000 658.500000 487.650000 ;
      RECT 616.500000 486.350000 649.500000 487.650000 ;
      RECT 607.500000 486.350000 608.500000 487.650000 ;
      RECT 566.500000 486.350000 599.500000 487.650000 ;
      RECT 557.500000 486.350000 558.500000 487.650000 ;
      RECT 516.500000 486.350000 549.500000 487.650000 ;
      RECT 507.500000 486.350000 508.500000 487.650000 ;
      RECT 466.500000 486.350000 499.500000 487.650000 ;
      RECT 457.500000 486.350000 458.500000 487.650000 ;
      RECT 416.500000 486.350000 449.500000 487.650000 ;
      RECT 407.500000 486.350000 408.500000 487.650000 ;
      RECT 382.500000 486.350000 399.500000 487.650000 ;
      RECT 366.500000 486.350000 369.500000 489.650000 ;
      RECT 357.500000 486.350000 358.500000 487.650000 ;
      RECT 316.500000 486.350000 349.500000 487.650000 ;
      RECT 307.500000 486.350000 308.500000 487.650000 ;
      RECT 266.500000 486.350000 299.500000 487.650000 ;
      RECT 257.500000 486.350000 258.500000 487.650000 ;
      RECT 216.500000 486.350000 249.500000 487.650000 ;
      RECT 207.500000 486.350000 208.500000 487.650000 ;
      RECT 166.500000 486.350000 199.500000 487.650000 ;
      RECT 157.500000 486.350000 158.500000 487.650000 ;
      RECT 116.500000 486.350000 149.500000 487.650000 ;
      RECT 107.500000 486.350000 108.500000 487.650000 ;
      RECT 66.500000 486.350000 99.500000 487.650000 ;
      RECT 57.500000 486.350000 58.500000 487.650000 ;
      RECT 29.500000 486.350000 49.500000 487.650000 ;
      RECT 15.500000 486.350000 16.500000 487.650000 ;
      RECT 1157.500000 485.650000 1183.980000 486.350000 ;
      RECT 707.500000 485.650000 733.500000 486.350000 ;
      RECT 657.500000 485.650000 699.500000 486.350000 ;
      RECT 607.500000 485.650000 649.500000 486.350000 ;
      RECT 557.500000 485.650000 599.500000 486.350000 ;
      RECT 507.500000 485.650000 549.500000 486.350000 ;
      RECT 457.500000 485.650000 499.500000 486.350000 ;
      RECT 407.500000 485.650000 449.500000 486.350000 ;
      RECT 357.500000 485.650000 399.500000 486.350000 ;
      RECT 307.500000 485.650000 349.500000 486.350000 ;
      RECT 257.500000 485.650000 299.500000 486.350000 ;
      RECT 207.500000 485.650000 249.500000 486.350000 ;
      RECT 157.500000 485.650000 199.500000 486.350000 ;
      RECT 107.500000 485.650000 149.500000 486.350000 ;
      RECT 57.500000 485.650000 99.500000 486.350000 ;
      RECT 15.500000 485.650000 49.500000 486.350000 ;
      RECT 1157.500000 484.350000 1158.500000 485.650000 ;
      RECT 1139.000000 484.350000 1149.500000 487.650000 ;
      RECT 746.500000 484.350000 749.000000 487.650000 ;
      RECT 732.500000 484.350000 733.500000 485.650000 ;
      RECT 707.500000 484.350000 708.500000 485.650000 ;
      RECT 666.500000 484.350000 699.500000 485.650000 ;
      RECT 657.500000 484.350000 658.500000 485.650000 ;
      RECT 616.500000 484.350000 649.500000 485.650000 ;
      RECT 607.500000 484.350000 608.500000 485.650000 ;
      RECT 566.500000 484.350000 599.500000 485.650000 ;
      RECT 557.500000 484.350000 558.500000 485.650000 ;
      RECT 516.500000 484.350000 549.500000 485.650000 ;
      RECT 507.500000 484.350000 508.500000 485.650000 ;
      RECT 466.500000 484.350000 499.500000 485.650000 ;
      RECT 457.500000 484.350000 458.500000 485.650000 ;
      RECT 416.500000 484.350000 449.500000 485.650000 ;
      RECT 407.500000 484.350000 408.500000 485.650000 ;
      RECT 382.500000 484.350000 399.500000 485.650000 ;
      RECT 357.500000 484.350000 358.500000 485.650000 ;
      RECT 316.500000 484.350000 349.500000 485.650000 ;
      RECT 307.500000 484.350000 308.500000 485.650000 ;
      RECT 266.500000 484.350000 299.500000 485.650000 ;
      RECT 257.500000 484.350000 258.500000 485.650000 ;
      RECT 216.500000 484.350000 249.500000 485.650000 ;
      RECT 207.500000 484.350000 208.500000 485.650000 ;
      RECT 166.500000 484.350000 199.500000 485.650000 ;
      RECT 157.500000 484.350000 158.500000 485.650000 ;
      RECT 116.500000 484.350000 149.500000 485.650000 ;
      RECT 107.500000 484.350000 108.500000 485.650000 ;
      RECT 66.500000 484.350000 99.500000 485.650000 ;
      RECT 57.500000 484.350000 58.500000 485.650000 ;
      RECT 29.500000 484.350000 49.500000 485.650000 ;
      RECT 15.500000 484.350000 16.500000 485.650000 ;
      RECT 2.020000 484.350000 2.500000 487.170000 ;
      RECT 2.020000 484.070000 16.500000 484.350000 ;
      RECT 1166.500000 484.065000 1183.980000 485.650000 ;
      RECT 1139.000000 483.650000 1158.500000 484.350000 ;
      RECT 732.500000 483.650000 749.000000 484.350000 ;
      RECT 666.500000 483.650000 708.500000 484.350000 ;
      RECT 616.500000 483.650000 658.500000 484.350000 ;
      RECT 566.500000 483.650000 608.500000 484.350000 ;
      RECT 516.500000 483.650000 558.500000 484.350000 ;
      RECT 466.500000 483.650000 508.500000 484.350000 ;
      RECT 416.500000 483.650000 458.500000 484.350000 ;
      RECT 382.500000 483.650000 408.500000 484.350000 ;
      RECT 316.500000 483.650000 358.500000 484.350000 ;
      RECT 266.500000 483.650000 308.500000 484.350000 ;
      RECT 216.500000 483.650000 258.500000 484.350000 ;
      RECT 166.500000 483.650000 208.500000 484.350000 ;
      RECT 116.500000 483.650000 158.500000 484.350000 ;
      RECT 66.500000 483.650000 108.500000 484.350000 ;
      RECT 29.500000 483.650000 58.500000 484.350000 ;
      RECT 0.000000 483.650000 16.500000 484.070000 ;
      RECT 1166.500000 482.350000 1186.000000 484.065000 ;
      RECT 1157.500000 482.350000 1158.500000 483.650000 ;
      RECT 732.500000 482.350000 733.500000 483.650000 ;
      RECT 716.500000 482.350000 719.500000 485.650000 ;
      RECT 707.500000 482.350000 708.500000 483.650000 ;
      RECT 666.500000 482.350000 699.500000 483.650000 ;
      RECT 657.500000 482.350000 658.500000 483.650000 ;
      RECT 616.500000 482.350000 649.500000 483.650000 ;
      RECT 607.500000 482.350000 608.500000 483.650000 ;
      RECT 566.500000 482.350000 599.500000 483.650000 ;
      RECT 557.500000 482.350000 558.500000 483.650000 ;
      RECT 516.500000 482.350000 549.500000 483.650000 ;
      RECT 507.500000 482.350000 508.500000 483.650000 ;
      RECT 466.500000 482.350000 499.500000 483.650000 ;
      RECT 457.500000 482.350000 458.500000 483.650000 ;
      RECT 416.500000 482.350000 449.500000 483.650000 ;
      RECT 407.500000 482.350000 408.500000 483.650000 ;
      RECT 382.500000 482.350000 399.500000 483.650000 ;
      RECT 366.500000 482.350000 369.500000 485.650000 ;
      RECT 357.500000 482.350000 358.500000 483.650000 ;
      RECT 316.500000 482.350000 349.500000 483.650000 ;
      RECT 307.500000 482.350000 308.500000 483.650000 ;
      RECT 266.500000 482.350000 299.500000 483.650000 ;
      RECT 257.500000 482.350000 258.500000 483.650000 ;
      RECT 216.500000 482.350000 249.500000 483.650000 ;
      RECT 207.500000 482.350000 208.500000 483.650000 ;
      RECT 166.500000 482.350000 199.500000 483.650000 ;
      RECT 157.500000 482.350000 158.500000 483.650000 ;
      RECT 116.500000 482.350000 149.500000 483.650000 ;
      RECT 107.500000 482.350000 108.500000 483.650000 ;
      RECT 66.500000 482.350000 99.500000 483.650000 ;
      RECT 57.500000 482.350000 58.500000 483.650000 ;
      RECT 29.500000 482.350000 49.500000 483.650000 ;
      RECT 15.500000 482.350000 16.500000 483.650000 ;
      RECT 1157.500000 481.650000 1186.000000 482.350000 ;
      RECT 707.500000 481.650000 733.500000 482.350000 ;
      RECT 657.500000 481.650000 699.500000 482.350000 ;
      RECT 607.500000 481.650000 649.500000 482.350000 ;
      RECT 557.500000 481.650000 599.500000 482.350000 ;
      RECT 507.500000 481.650000 549.500000 482.350000 ;
      RECT 457.500000 481.650000 499.500000 482.350000 ;
      RECT 407.500000 481.650000 449.500000 482.350000 ;
      RECT 357.500000 481.650000 399.500000 482.350000 ;
      RECT 307.500000 481.650000 349.500000 482.350000 ;
      RECT 257.500000 481.650000 299.500000 482.350000 ;
      RECT 207.500000 481.650000 249.500000 482.350000 ;
      RECT 157.500000 481.650000 199.500000 482.350000 ;
      RECT 107.500000 481.650000 149.500000 482.350000 ;
      RECT 57.500000 481.650000 99.500000 482.350000 ;
      RECT 15.500000 481.650000 49.500000 482.350000 ;
      RECT 1166.500000 481.485000 1186.000000 481.650000 ;
      RECT 1157.500000 480.350000 1158.500000 481.650000 ;
      RECT 1139.000000 480.350000 1149.500000 483.650000 ;
      RECT 746.500000 480.350000 749.000000 483.650000 ;
      RECT 732.500000 480.350000 733.500000 481.650000 ;
      RECT 707.500000 480.350000 708.500000 481.650000 ;
      RECT 666.500000 480.350000 699.500000 481.650000 ;
      RECT 657.500000 480.350000 658.500000 481.650000 ;
      RECT 616.500000 480.350000 649.500000 481.650000 ;
      RECT 607.500000 480.350000 608.500000 481.650000 ;
      RECT 566.500000 480.350000 599.500000 481.650000 ;
      RECT 557.500000 480.350000 558.500000 481.650000 ;
      RECT 516.500000 480.350000 549.500000 481.650000 ;
      RECT 507.500000 480.350000 508.500000 481.650000 ;
      RECT 466.500000 480.350000 499.500000 481.650000 ;
      RECT 457.500000 480.350000 458.500000 481.650000 ;
      RECT 416.500000 480.350000 449.500000 481.650000 ;
      RECT 407.500000 480.350000 408.500000 481.650000 ;
      RECT 382.500000 480.350000 399.500000 481.650000 ;
      RECT 357.500000 480.350000 358.500000 481.650000 ;
      RECT 316.500000 480.350000 349.500000 481.650000 ;
      RECT 307.500000 480.350000 308.500000 481.650000 ;
      RECT 266.500000 480.350000 299.500000 481.650000 ;
      RECT 257.500000 480.350000 258.500000 481.650000 ;
      RECT 216.500000 480.350000 249.500000 481.650000 ;
      RECT 207.500000 480.350000 208.500000 481.650000 ;
      RECT 166.500000 480.350000 199.500000 481.650000 ;
      RECT 157.500000 480.350000 158.500000 481.650000 ;
      RECT 116.500000 480.350000 149.500000 481.650000 ;
      RECT 107.500000 480.350000 108.500000 481.650000 ;
      RECT 66.500000 480.350000 99.500000 481.650000 ;
      RECT 57.500000 480.350000 58.500000 481.650000 ;
      RECT 29.500000 480.350000 49.500000 481.650000 ;
      RECT 15.500000 480.350000 16.500000 481.650000 ;
      RECT 0.000000 480.350000 2.500000 483.650000 ;
      RECT 1139.000000 479.650000 1158.500000 480.350000 ;
      RECT 732.500000 479.650000 749.000000 480.350000 ;
      RECT 666.500000 479.650000 708.500000 480.350000 ;
      RECT 616.500000 479.650000 658.500000 480.350000 ;
      RECT 566.500000 479.650000 608.500000 480.350000 ;
      RECT 516.500000 479.650000 558.500000 480.350000 ;
      RECT 466.500000 479.650000 508.500000 480.350000 ;
      RECT 416.500000 479.650000 458.500000 480.350000 ;
      RECT 382.500000 479.650000 408.500000 480.350000 ;
      RECT 316.500000 479.650000 358.500000 480.350000 ;
      RECT 266.500000 479.650000 308.500000 480.350000 ;
      RECT 216.500000 479.650000 258.500000 480.350000 ;
      RECT 166.500000 479.650000 208.500000 480.350000 ;
      RECT 116.500000 479.650000 158.500000 480.350000 ;
      RECT 66.500000 479.650000 108.500000 480.350000 ;
      RECT 29.500000 479.650000 58.500000 480.350000 ;
      RECT 0.000000 479.650000 16.500000 480.350000 ;
      RECT 1166.500000 478.385000 1183.980000 481.485000 ;
      RECT 1166.500000 478.350000 1186.000000 478.385000 ;
      RECT 1157.500000 478.350000 1158.500000 479.650000 ;
      RECT 732.500000 478.350000 733.500000 479.650000 ;
      RECT 716.500000 478.350000 719.500000 481.650000 ;
      RECT 707.500000 478.350000 708.500000 479.650000 ;
      RECT 666.500000 478.350000 699.500000 479.650000 ;
      RECT 657.500000 478.350000 658.500000 479.650000 ;
      RECT 616.500000 478.350000 649.500000 479.650000 ;
      RECT 607.500000 478.350000 608.500000 479.650000 ;
      RECT 566.500000 478.350000 599.500000 479.650000 ;
      RECT 557.500000 478.350000 558.500000 479.650000 ;
      RECT 516.500000 478.350000 549.500000 479.650000 ;
      RECT 507.500000 478.350000 508.500000 479.650000 ;
      RECT 466.500000 478.350000 499.500000 479.650000 ;
      RECT 457.500000 478.350000 458.500000 479.650000 ;
      RECT 416.500000 478.350000 449.500000 479.650000 ;
      RECT 407.500000 478.350000 408.500000 479.650000 ;
      RECT 382.500000 478.350000 399.500000 479.650000 ;
      RECT 366.500000 478.350000 369.500000 481.650000 ;
      RECT 357.500000 478.350000 358.500000 479.650000 ;
      RECT 316.500000 478.350000 349.500000 479.650000 ;
      RECT 307.500000 478.350000 308.500000 479.650000 ;
      RECT 266.500000 478.350000 299.500000 479.650000 ;
      RECT 257.500000 478.350000 258.500000 479.650000 ;
      RECT 216.500000 478.350000 249.500000 479.650000 ;
      RECT 207.500000 478.350000 208.500000 479.650000 ;
      RECT 166.500000 478.350000 199.500000 479.650000 ;
      RECT 157.500000 478.350000 158.500000 479.650000 ;
      RECT 116.500000 478.350000 149.500000 479.650000 ;
      RECT 107.500000 478.350000 108.500000 479.650000 ;
      RECT 66.500000 478.350000 99.500000 479.650000 ;
      RECT 57.500000 478.350000 58.500000 479.650000 ;
      RECT 29.500000 478.350000 49.500000 479.650000 ;
      RECT 15.500000 478.350000 16.500000 479.650000 ;
      RECT 1157.500000 477.650000 1186.000000 478.350000 ;
      RECT 707.500000 477.650000 733.500000 478.350000 ;
      RECT 657.500000 477.650000 699.500000 478.350000 ;
      RECT 607.500000 477.650000 649.500000 478.350000 ;
      RECT 557.500000 477.650000 599.500000 478.350000 ;
      RECT 507.500000 477.650000 549.500000 478.350000 ;
      RECT 457.500000 477.650000 499.500000 478.350000 ;
      RECT 407.500000 477.650000 449.500000 478.350000 ;
      RECT 357.500000 477.650000 399.500000 478.350000 ;
      RECT 307.500000 477.650000 349.500000 478.350000 ;
      RECT 257.500000 477.650000 299.500000 478.350000 ;
      RECT 207.500000 477.650000 249.500000 478.350000 ;
      RECT 157.500000 477.650000 199.500000 478.350000 ;
      RECT 107.500000 477.650000 149.500000 478.350000 ;
      RECT 57.500000 477.650000 99.500000 478.350000 ;
      RECT 15.500000 477.650000 49.500000 478.350000 ;
      RECT 1166.500000 477.525000 1186.000000 477.650000 ;
      RECT 0.000000 476.575000 2.500000 479.650000 ;
      RECT 1157.500000 476.350000 1158.500000 477.650000 ;
      RECT 1139.000000 476.350000 1149.500000 479.650000 ;
      RECT 746.500000 476.350000 749.000000 479.650000 ;
      RECT 732.500000 476.350000 733.500000 477.650000 ;
      RECT 707.500000 476.350000 708.500000 477.650000 ;
      RECT 666.500000 476.350000 699.500000 477.650000 ;
      RECT 657.500000 476.350000 658.500000 477.650000 ;
      RECT 616.500000 476.350000 649.500000 477.650000 ;
      RECT 607.500000 476.350000 608.500000 477.650000 ;
      RECT 566.500000 476.350000 599.500000 477.650000 ;
      RECT 557.500000 476.350000 558.500000 477.650000 ;
      RECT 516.500000 476.350000 549.500000 477.650000 ;
      RECT 507.500000 476.350000 508.500000 477.650000 ;
      RECT 466.500000 476.350000 499.500000 477.650000 ;
      RECT 457.500000 476.350000 458.500000 477.650000 ;
      RECT 416.500000 476.350000 449.500000 477.650000 ;
      RECT 407.500000 476.350000 408.500000 477.650000 ;
      RECT 366.500000 476.350000 399.500000 477.650000 ;
      RECT 357.500000 476.350000 358.500000 477.650000 ;
      RECT 316.500000 476.350000 349.500000 477.650000 ;
      RECT 307.500000 476.350000 308.500000 477.650000 ;
      RECT 266.500000 476.350000 299.500000 477.650000 ;
      RECT 257.500000 476.350000 258.500000 477.650000 ;
      RECT 216.500000 476.350000 249.500000 477.650000 ;
      RECT 207.500000 476.350000 208.500000 477.650000 ;
      RECT 166.500000 476.350000 199.500000 477.650000 ;
      RECT 157.500000 476.350000 158.500000 477.650000 ;
      RECT 116.500000 476.350000 149.500000 477.650000 ;
      RECT 107.500000 476.350000 108.500000 477.650000 ;
      RECT 66.500000 476.350000 99.500000 477.650000 ;
      RECT 57.500000 476.350000 58.500000 477.650000 ;
      RECT 29.500000 476.350000 49.500000 477.650000 ;
      RECT 15.500000 476.350000 16.500000 477.650000 ;
      RECT 2.020000 476.350000 2.500000 476.575000 ;
      RECT 1139.000000 475.650000 1158.500000 476.350000 ;
      RECT 732.500000 475.650000 749.000000 476.350000 ;
      RECT 666.500000 475.650000 708.500000 476.350000 ;
      RECT 616.500000 475.650000 658.500000 476.350000 ;
      RECT 566.500000 475.650000 608.500000 476.350000 ;
      RECT 516.500000 475.650000 558.500000 476.350000 ;
      RECT 466.500000 475.650000 508.500000 476.350000 ;
      RECT 416.500000 475.650000 458.500000 476.350000 ;
      RECT 366.500000 475.650000 408.500000 476.350000 ;
      RECT 316.500000 475.650000 358.500000 476.350000 ;
      RECT 266.500000 475.650000 308.500000 476.350000 ;
      RECT 216.500000 475.650000 258.500000 476.350000 ;
      RECT 166.500000 475.650000 208.500000 476.350000 ;
      RECT 116.500000 475.650000 158.500000 476.350000 ;
      RECT 66.500000 475.650000 108.500000 476.350000 ;
      RECT 29.500000 475.650000 58.500000 476.350000 ;
      RECT 2.020000 475.650000 16.500000 476.350000 ;
      RECT 1166.500000 474.425000 1183.980000 477.525000 ;
      RECT 1166.500000 474.350000 1186.000000 474.425000 ;
      RECT 1157.500000 474.350000 1158.500000 475.650000 ;
      RECT 732.500000 474.350000 733.500000 475.650000 ;
      RECT 716.500000 474.350000 719.500000 477.650000 ;
      RECT 707.500000 474.350000 708.500000 475.650000 ;
      RECT 666.500000 474.350000 699.500000 475.650000 ;
      RECT 657.500000 474.350000 658.500000 475.650000 ;
      RECT 616.500000 474.350000 649.500000 475.650000 ;
      RECT 607.500000 474.350000 608.500000 475.650000 ;
      RECT 566.500000 474.350000 599.500000 475.650000 ;
      RECT 557.500000 474.350000 558.500000 475.650000 ;
      RECT 516.500000 474.350000 549.500000 475.650000 ;
      RECT 507.500000 474.350000 508.500000 475.650000 ;
      RECT 466.500000 474.350000 499.500000 475.650000 ;
      RECT 457.500000 474.350000 458.500000 475.650000 ;
      RECT 416.500000 474.350000 449.500000 475.650000 ;
      RECT 407.500000 474.350000 408.500000 475.650000 ;
      RECT 366.500000 474.350000 399.500000 475.650000 ;
      RECT 357.500000 474.350000 358.500000 475.650000 ;
      RECT 316.500000 474.350000 349.500000 475.650000 ;
      RECT 307.500000 474.350000 308.500000 475.650000 ;
      RECT 266.500000 474.350000 299.500000 475.650000 ;
      RECT 257.500000 474.350000 258.500000 475.650000 ;
      RECT 216.500000 474.350000 249.500000 475.650000 ;
      RECT 207.500000 474.350000 208.500000 475.650000 ;
      RECT 166.500000 474.350000 199.500000 475.650000 ;
      RECT 157.500000 474.350000 158.500000 475.650000 ;
      RECT 116.500000 474.350000 149.500000 475.650000 ;
      RECT 107.500000 474.350000 108.500000 475.650000 ;
      RECT 66.500000 474.350000 99.500000 475.650000 ;
      RECT 57.500000 474.350000 58.500000 475.650000 ;
      RECT 29.500000 474.350000 49.500000 475.650000 ;
      RECT 15.500000 474.350000 16.500000 475.650000 ;
      RECT 1157.500000 473.650000 1186.000000 474.350000 ;
      RECT 707.500000 473.650000 733.500000 474.350000 ;
      RECT 657.500000 473.650000 699.500000 474.350000 ;
      RECT 607.500000 473.650000 649.500000 474.350000 ;
      RECT 557.500000 473.650000 599.500000 474.350000 ;
      RECT 507.500000 473.650000 549.500000 474.350000 ;
      RECT 457.500000 473.650000 499.500000 474.350000 ;
      RECT 407.500000 473.650000 449.500000 474.350000 ;
      RECT 357.500000 473.650000 399.500000 474.350000 ;
      RECT 307.500000 473.650000 349.500000 474.350000 ;
      RECT 257.500000 473.650000 299.500000 474.350000 ;
      RECT 207.500000 473.650000 249.500000 474.350000 ;
      RECT 157.500000 473.650000 199.500000 474.350000 ;
      RECT 107.500000 473.650000 149.500000 474.350000 ;
      RECT 57.500000 473.650000 99.500000 474.350000 ;
      RECT 15.500000 473.650000 49.500000 474.350000 ;
      RECT 2.020000 473.475000 2.500000 475.650000 ;
      RECT 0.000000 472.615000 2.500000 473.475000 ;
      RECT 1157.500000 472.350000 1158.500000 473.650000 ;
      RECT 1139.000000 472.350000 1149.500000 475.650000 ;
      RECT 746.500000 472.350000 749.000000 475.650000 ;
      RECT 732.500000 472.350000 733.500000 473.650000 ;
      RECT 707.500000 472.350000 708.500000 473.650000 ;
      RECT 666.500000 472.350000 699.500000 473.650000 ;
      RECT 657.500000 472.350000 658.500000 473.650000 ;
      RECT 616.500000 472.350000 649.500000 473.650000 ;
      RECT 607.500000 472.350000 608.500000 473.650000 ;
      RECT 566.500000 472.350000 599.500000 473.650000 ;
      RECT 557.500000 472.350000 558.500000 473.650000 ;
      RECT 516.500000 472.350000 549.500000 473.650000 ;
      RECT 507.500000 472.350000 508.500000 473.650000 ;
      RECT 466.500000 472.350000 499.500000 473.650000 ;
      RECT 457.500000 472.350000 458.500000 473.650000 ;
      RECT 416.500000 472.350000 449.500000 473.650000 ;
      RECT 407.500000 472.350000 408.500000 473.650000 ;
      RECT 366.500000 472.350000 399.500000 473.650000 ;
      RECT 357.500000 472.350000 358.500000 473.650000 ;
      RECT 316.500000 472.350000 349.500000 473.650000 ;
      RECT 307.500000 472.350000 308.500000 473.650000 ;
      RECT 266.500000 472.350000 299.500000 473.650000 ;
      RECT 257.500000 472.350000 258.500000 473.650000 ;
      RECT 216.500000 472.350000 249.500000 473.650000 ;
      RECT 207.500000 472.350000 208.500000 473.650000 ;
      RECT 166.500000 472.350000 199.500000 473.650000 ;
      RECT 157.500000 472.350000 158.500000 473.650000 ;
      RECT 116.500000 472.350000 149.500000 473.650000 ;
      RECT 107.500000 472.350000 108.500000 473.650000 ;
      RECT 66.500000 472.350000 99.500000 473.650000 ;
      RECT 57.500000 472.350000 58.500000 473.650000 ;
      RECT 29.500000 472.350000 49.500000 473.650000 ;
      RECT 15.500000 472.350000 16.500000 473.650000 ;
      RECT 2.020000 472.350000 2.500000 472.615000 ;
      RECT 1139.000000 471.650000 1158.500000 472.350000 ;
      RECT 732.500000 471.650000 749.000000 472.350000 ;
      RECT 666.500000 471.650000 708.500000 472.350000 ;
      RECT 616.500000 471.650000 658.500000 472.350000 ;
      RECT 566.500000 471.650000 608.500000 472.350000 ;
      RECT 516.500000 471.650000 558.500000 472.350000 ;
      RECT 466.500000 471.650000 508.500000 472.350000 ;
      RECT 416.500000 471.650000 458.500000 472.350000 ;
      RECT 366.500000 471.650000 408.500000 472.350000 ;
      RECT 316.500000 471.650000 358.500000 472.350000 ;
      RECT 266.500000 471.650000 308.500000 472.350000 ;
      RECT 216.500000 471.650000 258.500000 472.350000 ;
      RECT 166.500000 471.650000 208.500000 472.350000 ;
      RECT 116.500000 471.650000 158.500000 472.350000 ;
      RECT 66.500000 471.650000 108.500000 472.350000 ;
      RECT 29.500000 471.650000 58.500000 472.350000 ;
      RECT 2.020000 471.650000 16.500000 472.350000 ;
      RECT 1166.500000 470.350000 1186.000000 473.650000 ;
      RECT 1157.500000 470.350000 1158.500000 471.650000 ;
      RECT 732.500000 470.350000 733.500000 471.650000 ;
      RECT 716.500000 470.350000 719.500000 473.650000 ;
      RECT 707.500000 470.350000 708.500000 471.650000 ;
      RECT 666.500000 470.350000 699.500000 471.650000 ;
      RECT 657.500000 470.350000 658.500000 471.650000 ;
      RECT 616.500000 470.350000 649.500000 471.650000 ;
      RECT 607.500000 470.350000 608.500000 471.650000 ;
      RECT 566.500000 470.350000 599.500000 471.650000 ;
      RECT 557.500000 470.350000 558.500000 471.650000 ;
      RECT 516.500000 470.350000 549.500000 471.650000 ;
      RECT 507.500000 470.350000 508.500000 471.650000 ;
      RECT 466.500000 470.350000 499.500000 471.650000 ;
      RECT 457.500000 470.350000 458.500000 471.650000 ;
      RECT 416.500000 470.350000 449.500000 471.650000 ;
      RECT 407.500000 470.350000 408.500000 471.650000 ;
      RECT 366.500000 470.350000 399.500000 471.650000 ;
      RECT 357.500000 470.350000 358.500000 471.650000 ;
      RECT 316.500000 470.350000 349.500000 471.650000 ;
      RECT 307.500000 470.350000 308.500000 471.650000 ;
      RECT 266.500000 470.350000 299.500000 471.650000 ;
      RECT 257.500000 470.350000 258.500000 471.650000 ;
      RECT 216.500000 470.350000 249.500000 471.650000 ;
      RECT 207.500000 470.350000 208.500000 471.650000 ;
      RECT 166.500000 470.350000 199.500000 471.650000 ;
      RECT 157.500000 470.350000 158.500000 471.650000 ;
      RECT 116.500000 470.350000 149.500000 471.650000 ;
      RECT 107.500000 470.350000 108.500000 471.650000 ;
      RECT 66.500000 470.350000 99.500000 471.650000 ;
      RECT 57.500000 470.350000 58.500000 471.650000 ;
      RECT 29.500000 470.350000 49.500000 471.650000 ;
      RECT 15.500000 470.350000 16.500000 471.650000 ;
      RECT 1157.500000 469.650000 1186.000000 470.350000 ;
      RECT 707.500000 469.650000 733.500000 470.350000 ;
      RECT 657.500000 469.650000 699.500000 470.350000 ;
      RECT 607.500000 469.650000 649.500000 470.350000 ;
      RECT 557.500000 469.650000 599.500000 470.350000 ;
      RECT 507.500000 469.650000 549.500000 470.350000 ;
      RECT 457.500000 469.650000 499.500000 470.350000 ;
      RECT 407.500000 469.650000 449.500000 470.350000 ;
      RECT 357.500000 469.650000 399.500000 470.350000 ;
      RECT 307.500000 469.650000 349.500000 470.350000 ;
      RECT 257.500000 469.650000 299.500000 470.350000 ;
      RECT 207.500000 469.650000 249.500000 470.350000 ;
      RECT 157.500000 469.650000 199.500000 470.350000 ;
      RECT 107.500000 469.650000 149.500000 470.350000 ;
      RECT 57.500000 469.650000 99.500000 470.350000 ;
      RECT 15.500000 469.650000 49.500000 470.350000 ;
      RECT 2.020000 469.515000 2.500000 471.650000 ;
      RECT 1157.500000 468.350000 1158.500000 469.650000 ;
      RECT 1139.000000 468.350000 1149.500000 471.650000 ;
      RECT 746.500000 468.350000 749.000000 471.650000 ;
      RECT 732.500000 468.350000 733.500000 469.650000 ;
      RECT 707.500000 468.350000 708.500000 469.650000 ;
      RECT 666.500000 468.350000 699.500000 469.650000 ;
      RECT 657.500000 468.350000 658.500000 469.650000 ;
      RECT 616.500000 468.350000 649.500000 469.650000 ;
      RECT 607.500000 468.350000 608.500000 469.650000 ;
      RECT 566.500000 468.350000 599.500000 469.650000 ;
      RECT 557.500000 468.350000 558.500000 469.650000 ;
      RECT 516.500000 468.350000 549.500000 469.650000 ;
      RECT 507.500000 468.350000 508.500000 469.650000 ;
      RECT 466.500000 468.350000 499.500000 469.650000 ;
      RECT 457.500000 468.350000 458.500000 469.650000 ;
      RECT 416.500000 468.350000 449.500000 469.650000 ;
      RECT 407.500000 468.350000 408.500000 469.650000 ;
      RECT 366.500000 468.350000 399.500000 469.650000 ;
      RECT 357.500000 468.350000 358.500000 469.650000 ;
      RECT 316.500000 468.350000 349.500000 469.650000 ;
      RECT 307.500000 468.350000 308.500000 469.650000 ;
      RECT 266.500000 468.350000 299.500000 469.650000 ;
      RECT 257.500000 468.350000 258.500000 469.650000 ;
      RECT 216.500000 468.350000 249.500000 469.650000 ;
      RECT 207.500000 468.350000 208.500000 469.650000 ;
      RECT 166.500000 468.350000 199.500000 469.650000 ;
      RECT 157.500000 468.350000 158.500000 469.650000 ;
      RECT 116.500000 468.350000 149.500000 469.650000 ;
      RECT 107.500000 468.350000 108.500000 469.650000 ;
      RECT 66.500000 468.350000 99.500000 469.650000 ;
      RECT 57.500000 468.350000 58.500000 469.650000 ;
      RECT 29.500000 468.350000 49.500000 469.650000 ;
      RECT 15.500000 468.350000 16.500000 469.650000 ;
      RECT 0.000000 468.350000 2.500000 469.515000 ;
      RECT 1139.000000 467.650000 1158.500000 468.350000 ;
      RECT 732.500000 467.650000 749.000000 468.350000 ;
      RECT 666.500000 467.650000 708.500000 468.350000 ;
      RECT 616.500000 467.650000 658.500000 468.350000 ;
      RECT 566.500000 467.650000 608.500000 468.350000 ;
      RECT 516.500000 467.650000 558.500000 468.350000 ;
      RECT 466.500000 467.650000 508.500000 468.350000 ;
      RECT 416.500000 467.650000 458.500000 468.350000 ;
      RECT 366.500000 467.650000 408.500000 468.350000 ;
      RECT 316.500000 467.650000 358.500000 468.350000 ;
      RECT 266.500000 467.650000 308.500000 468.350000 ;
      RECT 216.500000 467.650000 258.500000 468.350000 ;
      RECT 166.500000 467.650000 208.500000 468.350000 ;
      RECT 116.500000 467.650000 158.500000 468.350000 ;
      RECT 66.500000 467.650000 108.500000 468.350000 ;
      RECT 29.500000 467.650000 58.500000 468.350000 ;
      RECT 0.000000 467.650000 16.500000 468.350000 ;
      RECT 0.000000 466.935000 2.500000 467.650000 ;
      RECT 1166.500000 466.930000 1186.000000 469.650000 ;
      RECT 1166.500000 466.350000 1183.980000 466.930000 ;
      RECT 1157.500000 466.350000 1158.500000 467.650000 ;
      RECT 732.500000 466.350000 733.500000 467.650000 ;
      RECT 716.500000 466.350000 719.500000 469.650000 ;
      RECT 707.500000 466.350000 708.500000 467.650000 ;
      RECT 666.500000 466.350000 699.500000 467.650000 ;
      RECT 657.500000 466.350000 658.500000 467.650000 ;
      RECT 616.500000 466.350000 649.500000 467.650000 ;
      RECT 607.500000 466.350000 608.500000 467.650000 ;
      RECT 566.500000 466.350000 599.500000 467.650000 ;
      RECT 557.500000 466.350000 558.500000 467.650000 ;
      RECT 516.500000 466.350000 549.500000 467.650000 ;
      RECT 507.500000 466.350000 508.500000 467.650000 ;
      RECT 466.500000 466.350000 499.500000 467.650000 ;
      RECT 457.500000 466.350000 458.500000 467.650000 ;
      RECT 416.500000 466.350000 449.500000 467.650000 ;
      RECT 407.500000 466.350000 408.500000 467.650000 ;
      RECT 366.500000 466.350000 399.500000 467.650000 ;
      RECT 357.500000 466.350000 358.500000 467.650000 ;
      RECT 316.500000 466.350000 349.500000 467.650000 ;
      RECT 307.500000 466.350000 308.500000 467.650000 ;
      RECT 266.500000 466.350000 299.500000 467.650000 ;
      RECT 257.500000 466.350000 258.500000 467.650000 ;
      RECT 216.500000 466.350000 249.500000 467.650000 ;
      RECT 207.500000 466.350000 208.500000 467.650000 ;
      RECT 166.500000 466.350000 199.500000 467.650000 ;
      RECT 157.500000 466.350000 158.500000 467.650000 ;
      RECT 116.500000 466.350000 149.500000 467.650000 ;
      RECT 107.500000 466.350000 108.500000 467.650000 ;
      RECT 66.500000 466.350000 99.500000 467.650000 ;
      RECT 57.500000 466.350000 58.500000 467.650000 ;
      RECT 29.500000 466.350000 49.500000 467.650000 ;
      RECT 15.500000 466.350000 16.500000 467.650000 ;
      RECT 1157.500000 465.650000 1183.980000 466.350000 ;
      RECT 707.500000 465.650000 733.500000 466.350000 ;
      RECT 657.500000 465.650000 699.500000 466.350000 ;
      RECT 607.500000 465.650000 649.500000 466.350000 ;
      RECT 557.500000 465.650000 599.500000 466.350000 ;
      RECT 507.500000 465.650000 549.500000 466.350000 ;
      RECT 457.500000 465.650000 499.500000 466.350000 ;
      RECT 407.500000 465.650000 449.500000 466.350000 ;
      RECT 357.500000 465.650000 399.500000 466.350000 ;
      RECT 307.500000 465.650000 349.500000 466.350000 ;
      RECT 257.500000 465.650000 299.500000 466.350000 ;
      RECT 207.500000 465.650000 249.500000 466.350000 ;
      RECT 157.500000 465.650000 199.500000 466.350000 ;
      RECT 107.500000 465.650000 149.500000 466.350000 ;
      RECT 57.500000 465.650000 99.500000 466.350000 ;
      RECT 15.500000 465.650000 49.500000 466.350000 ;
      RECT 1157.500000 464.350000 1158.500000 465.650000 ;
      RECT 1139.000000 464.350000 1149.500000 467.650000 ;
      RECT 746.500000 464.350000 749.000000 467.650000 ;
      RECT 732.500000 464.350000 733.500000 465.650000 ;
      RECT 707.500000 464.350000 708.500000 465.650000 ;
      RECT 666.500000 464.350000 699.500000 465.650000 ;
      RECT 657.500000 464.350000 658.500000 465.650000 ;
      RECT 616.500000 464.350000 649.500000 465.650000 ;
      RECT 607.500000 464.350000 608.500000 465.650000 ;
      RECT 566.500000 464.350000 599.500000 465.650000 ;
      RECT 557.500000 464.350000 558.500000 465.650000 ;
      RECT 516.500000 464.350000 549.500000 465.650000 ;
      RECT 507.500000 464.350000 508.500000 465.650000 ;
      RECT 466.500000 464.350000 499.500000 465.650000 ;
      RECT 457.500000 464.350000 458.500000 465.650000 ;
      RECT 416.500000 464.350000 449.500000 465.650000 ;
      RECT 407.500000 464.350000 408.500000 465.650000 ;
      RECT 366.500000 464.350000 399.500000 465.650000 ;
      RECT 357.500000 464.350000 358.500000 465.650000 ;
      RECT 316.500000 464.350000 349.500000 465.650000 ;
      RECT 307.500000 464.350000 308.500000 465.650000 ;
      RECT 266.500000 464.350000 299.500000 465.650000 ;
      RECT 257.500000 464.350000 258.500000 465.650000 ;
      RECT 216.500000 464.350000 249.500000 465.650000 ;
      RECT 207.500000 464.350000 208.500000 465.650000 ;
      RECT 166.500000 464.350000 199.500000 465.650000 ;
      RECT 157.500000 464.350000 158.500000 465.650000 ;
      RECT 116.500000 464.350000 149.500000 465.650000 ;
      RECT 107.500000 464.350000 108.500000 465.650000 ;
      RECT 66.500000 464.350000 99.500000 465.650000 ;
      RECT 57.500000 464.350000 58.500000 465.650000 ;
      RECT 29.500000 464.350000 49.500000 465.650000 ;
      RECT 15.500000 464.350000 16.500000 465.650000 ;
      RECT 2.020000 464.350000 2.500000 466.935000 ;
      RECT 2.020000 463.835000 16.500000 464.350000 ;
      RECT 1166.500000 463.830000 1183.980000 465.650000 ;
      RECT 1139.000000 463.650000 1158.500000 464.350000 ;
      RECT 732.500000 463.650000 749.000000 464.350000 ;
      RECT 666.500000 463.650000 708.500000 464.350000 ;
      RECT 616.500000 463.650000 658.500000 464.350000 ;
      RECT 566.500000 463.650000 608.500000 464.350000 ;
      RECT 516.500000 463.650000 558.500000 464.350000 ;
      RECT 466.500000 463.650000 508.500000 464.350000 ;
      RECT 416.500000 463.650000 458.500000 464.350000 ;
      RECT 366.500000 463.650000 408.500000 464.350000 ;
      RECT 316.500000 463.650000 358.500000 464.350000 ;
      RECT 266.500000 463.650000 308.500000 464.350000 ;
      RECT 216.500000 463.650000 258.500000 464.350000 ;
      RECT 166.500000 463.650000 208.500000 464.350000 ;
      RECT 116.500000 463.650000 158.500000 464.350000 ;
      RECT 66.500000 463.650000 108.500000 464.350000 ;
      RECT 29.500000 463.650000 58.500000 464.350000 ;
      RECT 0.000000 463.650000 16.500000 463.835000 ;
      RECT 1166.500000 462.350000 1186.000000 463.830000 ;
      RECT 1157.500000 462.350000 1158.500000 463.650000 ;
      RECT 732.500000 462.350000 733.500000 463.650000 ;
      RECT 716.500000 462.350000 719.500000 465.650000 ;
      RECT 707.500000 462.350000 708.500000 463.650000 ;
      RECT 666.500000 462.350000 699.500000 463.650000 ;
      RECT 657.500000 462.350000 658.500000 463.650000 ;
      RECT 616.500000 462.350000 649.500000 463.650000 ;
      RECT 607.500000 462.350000 608.500000 463.650000 ;
      RECT 566.500000 462.350000 599.500000 463.650000 ;
      RECT 557.500000 462.350000 558.500000 463.650000 ;
      RECT 516.500000 462.350000 549.500000 463.650000 ;
      RECT 507.500000 462.350000 508.500000 463.650000 ;
      RECT 466.500000 462.350000 499.500000 463.650000 ;
      RECT 457.500000 462.350000 458.500000 463.650000 ;
      RECT 416.500000 462.350000 449.500000 463.650000 ;
      RECT 407.500000 462.350000 408.500000 463.650000 ;
      RECT 366.500000 462.350000 399.500000 463.650000 ;
      RECT 357.500000 462.350000 358.500000 463.650000 ;
      RECT 316.500000 462.350000 349.500000 463.650000 ;
      RECT 307.500000 462.350000 308.500000 463.650000 ;
      RECT 266.500000 462.350000 299.500000 463.650000 ;
      RECT 257.500000 462.350000 258.500000 463.650000 ;
      RECT 216.500000 462.350000 249.500000 463.650000 ;
      RECT 207.500000 462.350000 208.500000 463.650000 ;
      RECT 166.500000 462.350000 199.500000 463.650000 ;
      RECT 157.500000 462.350000 158.500000 463.650000 ;
      RECT 116.500000 462.350000 149.500000 463.650000 ;
      RECT 107.500000 462.350000 108.500000 463.650000 ;
      RECT 66.500000 462.350000 99.500000 463.650000 ;
      RECT 57.500000 462.350000 58.500000 463.650000 ;
      RECT 29.500000 462.350000 49.500000 463.650000 ;
      RECT 15.500000 462.350000 16.500000 463.650000 ;
      RECT 1157.500000 461.650000 1186.000000 462.350000 ;
      RECT 707.500000 461.650000 733.500000 462.350000 ;
      RECT 657.500000 461.650000 699.500000 462.350000 ;
      RECT 607.500000 461.650000 649.500000 462.350000 ;
      RECT 557.500000 461.650000 599.500000 462.350000 ;
      RECT 507.500000 461.650000 549.500000 462.350000 ;
      RECT 457.500000 461.650000 499.500000 462.350000 ;
      RECT 407.500000 461.650000 449.500000 462.350000 ;
      RECT 357.500000 461.650000 399.500000 462.350000 ;
      RECT 307.500000 461.650000 349.500000 462.350000 ;
      RECT 207.500000 461.650000 249.500000 462.350000 ;
      RECT 107.500000 461.650000 149.500000 462.350000 ;
      RECT 57.500000 461.650000 99.500000 462.350000 ;
      RECT 15.500000 461.650000 49.500000 462.350000 ;
      RECT 1157.500000 460.350000 1158.500000 461.650000 ;
      RECT 1139.000000 460.350000 1149.500000 463.650000 ;
      RECT 746.500000 460.350000 749.000000 463.650000 ;
      RECT 732.500000 460.350000 733.500000 461.650000 ;
      RECT 707.500000 460.350000 708.500000 461.650000 ;
      RECT 666.500000 460.350000 699.500000 461.650000 ;
      RECT 657.500000 460.350000 658.500000 461.650000 ;
      RECT 616.500000 460.350000 649.500000 461.650000 ;
      RECT 607.500000 460.350000 608.500000 461.650000 ;
      RECT 566.500000 460.350000 599.500000 461.650000 ;
      RECT 557.500000 460.350000 558.500000 461.650000 ;
      RECT 516.500000 460.350000 549.500000 461.650000 ;
      RECT 507.500000 460.350000 508.500000 461.650000 ;
      RECT 466.500000 460.350000 499.500000 461.650000 ;
      RECT 457.500000 460.350000 458.500000 461.650000 ;
      RECT 416.500000 460.350000 449.500000 461.650000 ;
      RECT 407.500000 460.350000 408.500000 461.650000 ;
      RECT 366.500000 460.350000 399.500000 461.650000 ;
      RECT 357.500000 460.350000 358.500000 461.650000 ;
      RECT 316.500000 460.350000 349.500000 461.650000 ;
      RECT 307.500000 460.350000 308.500000 461.650000 ;
      RECT 257.500000 460.350000 299.500000 462.350000 ;
      RECT 216.500000 460.350000 249.500000 461.650000 ;
      RECT 207.500000 460.350000 208.500000 461.650000 ;
      RECT 157.500000 460.350000 199.500000 462.350000 ;
      RECT 116.500000 460.350000 149.500000 461.650000 ;
      RECT 107.500000 460.350000 108.500000 461.650000 ;
      RECT 66.500000 460.350000 99.500000 461.650000 ;
      RECT 57.500000 460.350000 58.500000 461.650000 ;
      RECT 29.500000 460.350000 49.500000 461.650000 ;
      RECT 15.500000 460.350000 16.500000 461.650000 ;
      RECT 0.000000 460.350000 2.500000 463.650000 ;
      RECT 1139.000000 459.650000 1158.500000 460.350000 ;
      RECT 732.500000 459.650000 749.000000 460.350000 ;
      RECT 666.500000 459.650000 708.500000 460.350000 ;
      RECT 616.500000 459.650000 658.500000 460.350000 ;
      RECT 566.500000 459.650000 608.500000 460.350000 ;
      RECT 516.500000 459.650000 558.500000 460.350000 ;
      RECT 466.500000 459.650000 508.500000 460.350000 ;
      RECT 416.500000 459.650000 458.500000 460.350000 ;
      RECT 366.500000 459.650000 408.500000 460.350000 ;
      RECT 316.500000 459.650000 358.500000 460.350000 ;
      RECT 216.500000 459.650000 308.500000 460.350000 ;
      RECT 116.500000 459.650000 208.500000 460.350000 ;
      RECT 66.500000 459.650000 108.500000 460.350000 ;
      RECT 29.500000 459.650000 58.500000 460.350000 ;
      RECT 0.000000 459.650000 16.500000 460.350000 ;
      RECT 1166.500000 458.350000 1186.000000 461.650000 ;
      RECT 1157.500000 458.350000 1158.500000 459.650000 ;
      RECT 732.500000 458.350000 733.500000 459.650000 ;
      RECT 716.500000 458.350000 719.500000 461.650000 ;
      RECT 707.500000 458.350000 708.500000 459.650000 ;
      RECT 666.500000 458.350000 699.500000 459.650000 ;
      RECT 657.500000 458.350000 658.500000 459.650000 ;
      RECT 616.500000 458.350000 649.500000 459.650000 ;
      RECT 607.500000 458.350000 608.500000 459.650000 ;
      RECT 566.500000 458.350000 599.500000 459.650000 ;
      RECT 557.500000 458.350000 558.500000 459.650000 ;
      RECT 516.500000 458.350000 549.500000 459.650000 ;
      RECT 507.500000 458.350000 508.500000 459.650000 ;
      RECT 466.500000 458.350000 499.500000 459.650000 ;
      RECT 457.500000 458.350000 458.500000 459.650000 ;
      RECT 416.500000 458.350000 449.500000 459.650000 ;
      RECT 407.500000 458.350000 408.500000 459.650000 ;
      RECT 366.500000 458.350000 399.500000 459.650000 ;
      RECT 357.500000 458.350000 358.500000 459.650000 ;
      RECT 316.500000 458.350000 349.500000 459.650000 ;
      RECT 307.500000 458.350000 308.500000 459.650000 ;
      RECT 216.500000 458.350000 249.500000 459.650000 ;
      RECT 207.500000 458.350000 208.500000 459.650000 ;
      RECT 116.500000 458.350000 149.500000 459.650000 ;
      RECT 107.500000 458.350000 108.500000 459.650000 ;
      RECT 66.500000 458.350000 99.500000 459.650000 ;
      RECT 57.500000 458.350000 58.500000 459.650000 ;
      RECT 29.500000 458.350000 49.500000 459.650000 ;
      RECT 15.500000 458.350000 16.500000 459.650000 ;
      RECT 1157.500000 457.650000 1186.000000 458.350000 ;
      RECT 707.500000 457.650000 733.500000 458.350000 ;
      RECT 657.500000 457.650000 699.500000 458.350000 ;
      RECT 607.500000 457.650000 649.500000 458.350000 ;
      RECT 557.500000 457.650000 599.500000 458.350000 ;
      RECT 507.500000 457.650000 549.500000 458.350000 ;
      RECT 457.500000 457.650000 499.500000 458.350000 ;
      RECT 407.500000 457.650000 449.500000 458.350000 ;
      RECT 357.500000 457.650000 399.500000 458.350000 ;
      RECT 307.500000 457.650000 349.500000 458.350000 ;
      RECT 207.500000 457.650000 249.500000 458.350000 ;
      RECT 107.500000 457.650000 149.500000 458.350000 ;
      RECT 57.500000 457.650000 99.500000 458.350000 ;
      RECT 15.500000 457.650000 49.500000 458.350000 ;
      RECT 1157.500000 456.350000 1158.500000 457.650000 ;
      RECT 1139.000000 456.350000 1149.500000 459.650000 ;
      RECT 746.500000 456.350000 749.000000 459.650000 ;
      RECT 732.500000 456.350000 733.500000 457.650000 ;
      RECT 707.500000 456.350000 708.500000 457.650000 ;
      RECT 666.500000 456.350000 699.500000 457.650000 ;
      RECT 657.500000 456.350000 658.500000 457.650000 ;
      RECT 616.500000 456.350000 649.500000 457.650000 ;
      RECT 607.500000 456.350000 608.500000 457.650000 ;
      RECT 566.500000 456.350000 599.500000 457.650000 ;
      RECT 557.500000 456.350000 558.500000 457.650000 ;
      RECT 516.500000 456.350000 549.500000 457.650000 ;
      RECT 507.500000 456.350000 508.500000 457.650000 ;
      RECT 466.500000 456.350000 499.500000 457.650000 ;
      RECT 457.500000 456.350000 458.500000 457.650000 ;
      RECT 416.500000 456.350000 449.500000 457.650000 ;
      RECT 407.500000 456.350000 408.500000 457.650000 ;
      RECT 366.500000 456.350000 399.500000 457.650000 ;
      RECT 357.500000 456.350000 358.500000 457.650000 ;
      RECT 316.500000 456.350000 349.500000 457.650000 ;
      RECT 307.500000 456.350000 308.500000 457.650000 ;
      RECT 257.500000 456.350000 299.500000 459.650000 ;
      RECT 216.500000 456.350000 249.500000 457.650000 ;
      RECT 207.500000 456.350000 208.500000 457.650000 ;
      RECT 157.500000 456.350000 199.500000 459.650000 ;
      RECT 116.500000 456.350000 149.500000 457.650000 ;
      RECT 107.500000 456.350000 108.500000 457.650000 ;
      RECT 66.500000 456.350000 99.500000 457.650000 ;
      RECT 57.500000 456.350000 58.500000 457.650000 ;
      RECT 29.500000 456.350000 49.500000 457.650000 ;
      RECT 15.500000 456.350000 16.500000 457.650000 ;
      RECT 0.000000 456.350000 2.500000 459.650000 ;
      RECT 1139.000000 455.650000 1158.500000 456.350000 ;
      RECT 732.500000 455.650000 749.000000 456.350000 ;
      RECT 666.500000 455.650000 708.500000 456.350000 ;
      RECT 616.500000 455.650000 658.500000 456.350000 ;
      RECT 566.500000 455.650000 608.500000 456.350000 ;
      RECT 516.500000 455.650000 558.500000 456.350000 ;
      RECT 466.500000 455.650000 508.500000 456.350000 ;
      RECT 416.500000 455.650000 458.500000 456.350000 ;
      RECT 366.500000 455.650000 408.500000 456.350000 ;
      RECT 316.500000 455.650000 358.500000 456.350000 ;
      RECT 216.500000 455.650000 308.500000 456.350000 ;
      RECT 116.500000 455.650000 208.500000 456.350000 ;
      RECT 66.500000 455.650000 108.500000 456.350000 ;
      RECT 29.500000 455.650000 58.500000 456.350000 ;
      RECT 0.000000 455.650000 16.500000 456.350000 ;
      RECT 1166.500000 454.350000 1186.000000 457.650000 ;
      RECT 1157.500000 454.350000 1158.500000 455.650000 ;
      RECT 732.500000 454.350000 733.500000 455.650000 ;
      RECT 716.500000 454.350000 719.500000 457.650000 ;
      RECT 707.500000 454.350000 708.500000 455.650000 ;
      RECT 666.500000 454.350000 699.500000 455.650000 ;
      RECT 657.500000 454.350000 658.500000 455.650000 ;
      RECT 616.500000 454.350000 649.500000 455.650000 ;
      RECT 607.500000 454.350000 608.500000 455.650000 ;
      RECT 566.500000 454.350000 599.500000 455.650000 ;
      RECT 557.500000 454.350000 558.500000 455.650000 ;
      RECT 516.500000 454.350000 549.500000 455.650000 ;
      RECT 507.500000 454.350000 508.500000 455.650000 ;
      RECT 466.500000 454.350000 499.500000 455.650000 ;
      RECT 457.500000 454.350000 458.500000 455.650000 ;
      RECT 416.500000 454.350000 449.500000 455.650000 ;
      RECT 407.500000 454.350000 408.500000 455.650000 ;
      RECT 366.500000 454.350000 399.500000 455.650000 ;
      RECT 357.500000 454.350000 358.500000 455.650000 ;
      RECT 316.500000 454.350000 349.500000 455.650000 ;
      RECT 307.500000 454.350000 308.500000 455.650000 ;
      RECT 216.500000 454.350000 249.500000 455.650000 ;
      RECT 207.500000 454.350000 208.500000 455.650000 ;
      RECT 116.500000 454.350000 149.500000 455.650000 ;
      RECT 107.500000 454.350000 108.500000 455.650000 ;
      RECT 66.500000 454.350000 99.500000 455.650000 ;
      RECT 57.500000 454.350000 58.500000 455.650000 ;
      RECT 29.500000 454.350000 49.500000 455.650000 ;
      RECT 15.500000 454.350000 16.500000 455.650000 ;
      RECT 1157.500000 453.650000 1186.000000 454.350000 ;
      RECT 707.500000 453.650000 733.500000 454.350000 ;
      RECT 657.500000 453.650000 699.500000 454.350000 ;
      RECT 607.500000 453.650000 649.500000 454.350000 ;
      RECT 557.500000 453.650000 599.500000 454.350000 ;
      RECT 507.500000 453.650000 549.500000 454.350000 ;
      RECT 457.500000 453.650000 499.500000 454.350000 ;
      RECT 407.500000 453.650000 449.500000 454.350000 ;
      RECT 357.500000 453.650000 399.500000 454.350000 ;
      RECT 307.500000 453.650000 349.500000 454.350000 ;
      RECT 207.500000 453.650000 249.500000 454.350000 ;
      RECT 107.500000 453.650000 149.500000 454.350000 ;
      RECT 57.500000 453.650000 99.500000 454.350000 ;
      RECT 15.500000 453.650000 49.500000 454.350000 ;
      RECT 1157.500000 452.350000 1158.500000 453.650000 ;
      RECT 1139.000000 452.350000 1149.500000 455.650000 ;
      RECT 746.500000 452.350000 749.000000 455.650000 ;
      RECT 732.500000 452.350000 733.500000 453.650000 ;
      RECT 707.500000 452.350000 708.500000 453.650000 ;
      RECT 666.500000 452.350000 699.500000 453.650000 ;
      RECT 657.500000 452.350000 658.500000 453.650000 ;
      RECT 616.500000 452.350000 649.500000 453.650000 ;
      RECT 607.500000 452.350000 608.500000 453.650000 ;
      RECT 566.500000 452.350000 599.500000 453.650000 ;
      RECT 557.500000 452.350000 558.500000 453.650000 ;
      RECT 516.500000 452.350000 549.500000 453.650000 ;
      RECT 507.500000 452.350000 508.500000 453.650000 ;
      RECT 466.500000 452.350000 499.500000 453.650000 ;
      RECT 457.500000 452.350000 458.500000 453.650000 ;
      RECT 416.500000 452.350000 449.500000 453.650000 ;
      RECT 407.500000 452.350000 408.500000 453.650000 ;
      RECT 366.500000 452.350000 399.500000 453.650000 ;
      RECT 357.500000 452.350000 358.500000 453.650000 ;
      RECT 316.500000 452.350000 349.500000 453.650000 ;
      RECT 307.500000 452.350000 308.500000 453.650000 ;
      RECT 257.500000 452.350000 299.500000 455.650000 ;
      RECT 216.500000 452.350000 249.500000 453.650000 ;
      RECT 207.500000 452.350000 208.500000 453.650000 ;
      RECT 157.500000 452.350000 199.500000 455.650000 ;
      RECT 116.500000 452.350000 149.500000 453.650000 ;
      RECT 107.500000 452.350000 108.500000 453.650000 ;
      RECT 66.500000 452.350000 99.500000 453.650000 ;
      RECT 57.500000 452.350000 58.500000 453.650000 ;
      RECT 29.500000 452.350000 49.500000 453.650000 ;
      RECT 15.500000 452.350000 16.500000 453.650000 ;
      RECT 0.000000 452.350000 2.500000 455.650000 ;
      RECT 1139.000000 451.650000 1158.500000 452.350000 ;
      RECT 732.500000 451.650000 749.000000 452.350000 ;
      RECT 666.500000 451.650000 708.500000 452.350000 ;
      RECT 616.500000 451.650000 658.500000 452.350000 ;
      RECT 566.500000 451.650000 608.500000 452.350000 ;
      RECT 516.500000 451.650000 558.500000 452.350000 ;
      RECT 466.500000 451.650000 508.500000 452.350000 ;
      RECT 416.500000 451.650000 458.500000 452.350000 ;
      RECT 366.500000 451.650000 408.500000 452.350000 ;
      RECT 316.500000 451.650000 358.500000 452.350000 ;
      RECT 216.500000 451.650000 308.500000 452.350000 ;
      RECT 116.500000 451.650000 208.500000 452.350000 ;
      RECT 66.500000 451.650000 108.500000 452.350000 ;
      RECT 29.500000 451.650000 58.500000 452.350000 ;
      RECT 0.000000 451.650000 16.500000 452.350000 ;
      RECT 1166.500000 450.350000 1186.000000 453.650000 ;
      RECT 1157.500000 450.350000 1158.500000 451.650000 ;
      RECT 732.500000 450.350000 733.500000 451.650000 ;
      RECT 716.500000 450.350000 719.500000 453.650000 ;
      RECT 707.500000 450.350000 708.500000 451.650000 ;
      RECT 666.500000 450.350000 699.500000 451.650000 ;
      RECT 657.500000 450.350000 658.500000 451.650000 ;
      RECT 616.500000 450.350000 649.500000 451.650000 ;
      RECT 607.500000 450.350000 608.500000 451.650000 ;
      RECT 566.500000 450.350000 599.500000 451.650000 ;
      RECT 557.500000 450.350000 558.500000 451.650000 ;
      RECT 516.500000 450.350000 549.500000 451.650000 ;
      RECT 507.500000 450.350000 508.500000 451.650000 ;
      RECT 466.500000 450.350000 499.500000 451.650000 ;
      RECT 457.500000 450.350000 458.500000 451.650000 ;
      RECT 416.500000 450.350000 449.500000 451.650000 ;
      RECT 407.500000 450.350000 408.500000 451.650000 ;
      RECT 366.500000 450.350000 399.500000 451.650000 ;
      RECT 357.500000 450.350000 358.500000 451.650000 ;
      RECT 316.500000 450.350000 349.500000 451.650000 ;
      RECT 307.500000 450.350000 308.500000 451.650000 ;
      RECT 216.500000 450.350000 299.500000 451.650000 ;
      RECT 207.500000 450.350000 208.500000 451.650000 ;
      RECT 116.500000 450.350000 199.500000 451.650000 ;
      RECT 107.500000 450.350000 108.500000 451.650000 ;
      RECT 66.500000 450.350000 99.500000 451.650000 ;
      RECT 57.500000 450.350000 58.500000 451.650000 ;
      RECT 29.500000 450.350000 49.500000 451.650000 ;
      RECT 15.500000 450.350000 16.500000 451.650000 ;
      RECT 1157.500000 449.650000 1186.000000 450.350000 ;
      RECT 707.500000 449.650000 733.500000 450.350000 ;
      RECT 657.500000 449.650000 699.500000 450.350000 ;
      RECT 607.500000 449.650000 649.500000 450.350000 ;
      RECT 557.500000 449.650000 599.500000 450.350000 ;
      RECT 507.500000 449.650000 549.500000 450.350000 ;
      RECT 457.500000 449.650000 499.500000 450.350000 ;
      RECT 407.500000 449.650000 449.500000 450.350000 ;
      RECT 357.500000 449.650000 399.500000 450.350000 ;
      RECT 307.500000 449.650000 349.500000 450.350000 ;
      RECT 207.500000 449.650000 299.500000 450.350000 ;
      RECT 107.500000 449.650000 199.500000 450.350000 ;
      RECT 57.500000 449.650000 99.500000 450.350000 ;
      RECT 15.500000 449.650000 49.500000 450.350000 ;
      RECT 1157.500000 448.350000 1158.500000 449.650000 ;
      RECT 1139.000000 448.350000 1149.500000 451.650000 ;
      RECT 746.500000 448.350000 749.000000 451.650000 ;
      RECT 732.500000 448.350000 733.500000 449.650000 ;
      RECT 707.500000 448.350000 708.500000 449.650000 ;
      RECT 666.500000 448.350000 699.500000 449.650000 ;
      RECT 657.500000 448.350000 658.500000 449.650000 ;
      RECT 616.500000 448.350000 649.500000 449.650000 ;
      RECT 607.500000 448.350000 608.500000 449.650000 ;
      RECT 566.500000 448.350000 599.500000 449.650000 ;
      RECT 557.500000 448.350000 558.500000 449.650000 ;
      RECT 516.500000 448.350000 549.500000 449.650000 ;
      RECT 507.500000 448.350000 508.500000 449.650000 ;
      RECT 466.500000 448.350000 499.500000 449.650000 ;
      RECT 457.500000 448.350000 458.500000 449.650000 ;
      RECT 416.500000 448.350000 449.500000 449.650000 ;
      RECT 407.500000 448.350000 408.500000 449.650000 ;
      RECT 366.500000 448.350000 399.500000 449.650000 ;
      RECT 357.500000 448.350000 358.500000 449.650000 ;
      RECT 316.500000 448.350000 349.500000 449.650000 ;
      RECT 307.500000 448.350000 308.500000 449.650000 ;
      RECT 216.500000 448.350000 299.500000 449.650000 ;
      RECT 207.500000 448.350000 208.500000 449.650000 ;
      RECT 116.500000 448.350000 199.500000 449.650000 ;
      RECT 107.500000 448.350000 108.500000 449.650000 ;
      RECT 66.500000 448.350000 99.500000 449.650000 ;
      RECT 57.500000 448.350000 58.500000 449.650000 ;
      RECT 29.500000 448.350000 49.500000 449.650000 ;
      RECT 15.500000 448.350000 16.500000 449.650000 ;
      RECT 0.000000 448.350000 2.500000 451.650000 ;
      RECT 1139.000000 447.650000 1158.500000 448.350000 ;
      RECT 732.500000 447.650000 749.000000 448.350000 ;
      RECT 666.500000 447.650000 708.500000 448.350000 ;
      RECT 616.500000 447.650000 658.500000 448.350000 ;
      RECT 566.500000 447.650000 608.500000 448.350000 ;
      RECT 516.500000 447.650000 558.500000 448.350000 ;
      RECT 466.500000 447.650000 508.500000 448.350000 ;
      RECT 416.500000 447.650000 458.500000 448.350000 ;
      RECT 366.500000 447.650000 408.500000 448.350000 ;
      RECT 316.500000 447.650000 358.500000 448.350000 ;
      RECT 216.500000 447.650000 308.500000 448.350000 ;
      RECT 116.500000 447.650000 208.500000 448.350000 ;
      RECT 66.500000 447.650000 108.500000 448.350000 ;
      RECT 29.500000 447.650000 58.500000 448.350000 ;
      RECT 0.000000 447.650000 16.500000 448.350000 ;
      RECT 1166.500000 446.350000 1186.000000 449.650000 ;
      RECT 1157.500000 446.350000 1158.500000 447.650000 ;
      RECT 732.500000 446.350000 733.500000 447.650000 ;
      RECT 716.500000 446.350000 719.500000 449.650000 ;
      RECT 707.500000 446.350000 708.500000 447.650000 ;
      RECT 666.500000 446.350000 699.500000 447.650000 ;
      RECT 657.500000 446.350000 658.500000 447.650000 ;
      RECT 616.500000 446.350000 649.500000 447.650000 ;
      RECT 607.500000 446.350000 608.500000 447.650000 ;
      RECT 566.500000 446.350000 599.500000 447.650000 ;
      RECT 557.500000 446.350000 558.500000 447.650000 ;
      RECT 516.500000 446.350000 549.500000 447.650000 ;
      RECT 507.500000 446.350000 508.500000 447.650000 ;
      RECT 466.500000 446.350000 499.500000 447.650000 ;
      RECT 457.500000 446.350000 458.500000 447.650000 ;
      RECT 416.500000 446.350000 449.500000 447.650000 ;
      RECT 407.500000 446.350000 408.500000 447.650000 ;
      RECT 366.500000 446.350000 399.500000 447.650000 ;
      RECT 357.500000 446.350000 358.500000 447.650000 ;
      RECT 316.500000 446.350000 349.500000 447.650000 ;
      RECT 307.500000 446.350000 308.500000 447.650000 ;
      RECT 216.500000 446.350000 299.500000 447.650000 ;
      RECT 207.500000 446.350000 208.500000 447.650000 ;
      RECT 116.500000 446.350000 199.500000 447.650000 ;
      RECT 107.500000 446.350000 108.500000 447.650000 ;
      RECT 66.500000 446.350000 99.500000 447.650000 ;
      RECT 57.500000 446.350000 58.500000 447.650000 ;
      RECT 29.500000 446.350000 49.500000 447.650000 ;
      RECT 15.500000 446.350000 16.500000 447.650000 ;
      RECT 1139.000000 446.000000 1149.500000 447.650000 ;
      RECT 746.500000 446.000000 749.000000 447.650000 ;
      RECT 1157.500000 445.650000 1186.000000 446.350000 ;
      RECT 1055.460000 445.650000 1149.500000 446.000000 ;
      RECT 1009.630000 445.650000 1019.115000 446.000000 ;
      RECT 886.205000 445.650000 1006.530000 446.000000 ;
      RECT 746.500000 445.650000 878.305000 446.000000 ;
      RECT 707.500000 445.650000 733.500000 446.350000 ;
      RECT 657.500000 445.650000 699.500000 446.350000 ;
      RECT 607.500000 445.650000 649.500000 446.350000 ;
      RECT 557.500000 445.650000 599.500000 446.350000 ;
      RECT 507.500000 445.650000 549.500000 446.350000 ;
      RECT 457.500000 445.650000 499.500000 446.350000 ;
      RECT 407.500000 445.650000 449.500000 446.350000 ;
      RECT 357.500000 445.650000 399.500000 446.350000 ;
      RECT 307.500000 445.650000 349.500000 446.350000 ;
      RECT 207.500000 445.650000 299.500000 446.350000 ;
      RECT 107.500000 445.650000 199.500000 446.350000 ;
      RECT 57.500000 445.650000 99.500000 446.350000 ;
      RECT 15.500000 445.650000 49.500000 446.350000 ;
      RECT 1157.500000 444.350000 1158.500000 445.650000 ;
      RECT 1116.500000 444.350000 1149.500000 445.650000 ;
      RECT 746.500000 444.350000 758.500000 445.650000 ;
      RECT 732.500000 444.350000 733.500000 445.650000 ;
      RECT 707.500000 444.350000 708.500000 445.650000 ;
      RECT 666.500000 444.350000 699.500000 445.650000 ;
      RECT 657.500000 444.350000 658.500000 445.650000 ;
      RECT 616.500000 444.350000 649.500000 445.650000 ;
      RECT 607.500000 444.350000 608.500000 445.650000 ;
      RECT 566.500000 444.350000 599.500000 445.650000 ;
      RECT 557.500000 444.350000 558.500000 445.650000 ;
      RECT 516.500000 444.350000 549.500000 445.650000 ;
      RECT 507.500000 444.350000 508.500000 445.650000 ;
      RECT 466.500000 444.350000 499.500000 445.650000 ;
      RECT 457.500000 444.350000 458.500000 445.650000 ;
      RECT 416.500000 444.350000 449.500000 445.650000 ;
      RECT 407.500000 444.350000 408.500000 445.650000 ;
      RECT 366.500000 444.350000 399.500000 445.650000 ;
      RECT 357.500000 444.350000 358.500000 445.650000 ;
      RECT 316.500000 444.350000 349.500000 445.650000 ;
      RECT 307.500000 444.350000 308.500000 445.650000 ;
      RECT 216.500000 444.350000 299.500000 445.650000 ;
      RECT 207.500000 444.350000 208.500000 445.650000 ;
      RECT 116.500000 444.350000 199.500000 445.650000 ;
      RECT 107.500000 444.350000 108.500000 445.650000 ;
      RECT 66.500000 444.350000 99.500000 445.650000 ;
      RECT 57.500000 444.350000 58.500000 445.650000 ;
      RECT 29.500000 444.350000 49.500000 445.650000 ;
      RECT 15.500000 444.350000 16.500000 445.650000 ;
      RECT 0.000000 444.350000 2.500000 447.650000 ;
      RECT 1055.460000 443.980000 1058.500000 445.650000 ;
      RECT 1016.500000 443.980000 1019.115000 445.650000 ;
      RECT 966.500000 443.980000 1006.530000 445.650000 ;
      RECT 886.205000 443.980000 908.500000 445.650000 ;
      RECT 866.500000 443.980000 878.305000 445.650000 ;
      RECT 1166.500000 443.650000 1186.000000 445.650000 ;
      RECT 1116.500000 443.650000 1158.500000 444.350000 ;
      RECT 1066.500000 443.650000 1108.500000 445.650000 ;
      RECT 1016.500000 443.650000 1058.500000 443.980000 ;
      RECT 966.500000 443.650000 1008.500000 443.980000 ;
      RECT 916.500000 443.650000 958.500000 445.650000 ;
      RECT 866.500000 443.650000 908.500000 443.980000 ;
      RECT 816.500000 443.650000 858.500000 445.650000 ;
      RECT 766.500000 443.650000 808.500000 445.650000 ;
      RECT 732.500000 443.650000 758.500000 444.350000 ;
      RECT 666.500000 443.650000 708.500000 444.350000 ;
      RECT 616.500000 443.650000 658.500000 444.350000 ;
      RECT 566.500000 443.650000 608.500000 444.350000 ;
      RECT 516.500000 443.650000 558.500000 444.350000 ;
      RECT 466.500000 443.650000 508.500000 444.350000 ;
      RECT 416.500000 443.650000 458.500000 444.350000 ;
      RECT 366.500000 443.650000 408.500000 444.350000 ;
      RECT 316.500000 443.650000 358.500000 444.350000 ;
      RECT 216.500000 443.650000 308.500000 444.350000 ;
      RECT 116.500000 443.650000 208.500000 444.350000 ;
      RECT 66.500000 443.650000 108.500000 444.350000 ;
      RECT 29.500000 443.650000 58.500000 444.350000 ;
      RECT 0.000000 443.650000 16.500000 444.350000 ;
      RECT 1166.500000 442.350000 1170.500000 443.650000 ;
      RECT 1157.500000 442.350000 1158.500000 443.650000 ;
      RECT 1116.500000 442.350000 1149.500000 443.650000 ;
      RECT 1107.500000 442.350000 1108.500000 443.650000 ;
      RECT 1066.500000 442.350000 1099.500000 443.650000 ;
      RECT 1057.500000 442.350000 1058.500000 443.650000 ;
      RECT 1016.500000 442.350000 1049.500000 443.650000 ;
      RECT 1007.500000 442.350000 1008.500000 443.650000 ;
      RECT 966.500000 442.350000 999.500000 443.650000 ;
      RECT 957.500000 442.350000 958.500000 443.650000 ;
      RECT 916.500000 442.350000 949.500000 443.650000 ;
      RECT 907.500000 442.350000 908.500000 443.650000 ;
      RECT 866.500000 442.350000 899.500000 443.650000 ;
      RECT 857.500000 442.350000 858.500000 443.650000 ;
      RECT 816.500000 442.350000 849.500000 443.650000 ;
      RECT 807.500000 442.350000 808.500000 443.650000 ;
      RECT 766.500000 442.350000 799.500000 443.650000 ;
      RECT 757.500000 442.350000 758.500000 443.650000 ;
      RECT 732.500000 442.350000 733.500000 443.650000 ;
      RECT 716.500000 442.350000 719.500000 445.650000 ;
      RECT 707.500000 442.350000 708.500000 443.650000 ;
      RECT 666.500000 442.350000 699.500000 443.650000 ;
      RECT 657.500000 442.350000 658.500000 443.650000 ;
      RECT 616.500000 442.350000 649.500000 443.650000 ;
      RECT 607.500000 442.350000 608.500000 443.650000 ;
      RECT 566.500000 442.350000 599.500000 443.650000 ;
      RECT 557.500000 442.350000 558.500000 443.650000 ;
      RECT 516.500000 442.350000 549.500000 443.650000 ;
      RECT 507.500000 442.350000 508.500000 443.650000 ;
      RECT 466.500000 442.350000 499.500000 443.650000 ;
      RECT 457.500000 442.350000 458.500000 443.650000 ;
      RECT 416.500000 442.350000 449.500000 443.650000 ;
      RECT 407.500000 442.350000 408.500000 443.650000 ;
      RECT 366.500000 442.350000 399.500000 443.650000 ;
      RECT 357.500000 442.350000 358.500000 443.650000 ;
      RECT 316.500000 442.350000 349.500000 443.650000 ;
      RECT 307.500000 442.350000 308.500000 443.650000 ;
      RECT 216.500000 442.350000 299.500000 443.650000 ;
      RECT 207.500000 442.350000 208.500000 443.650000 ;
      RECT 116.500000 442.350000 199.500000 443.650000 ;
      RECT 107.500000 442.350000 108.500000 443.650000 ;
      RECT 66.500000 442.350000 99.500000 443.650000 ;
      RECT 57.500000 442.350000 58.500000 443.650000 ;
      RECT 29.500000 442.350000 49.500000 443.650000 ;
      RECT 15.500000 442.350000 16.500000 443.650000 ;
      RECT 1157.500000 441.650000 1170.500000 442.350000 ;
      RECT 1107.500000 441.650000 1149.500000 442.350000 ;
      RECT 1057.500000 441.650000 1099.500000 442.350000 ;
      RECT 1007.500000 441.650000 1049.500000 442.350000 ;
      RECT 957.500000 441.650000 999.500000 442.350000 ;
      RECT 907.500000 441.650000 949.500000 442.350000 ;
      RECT 857.500000 441.650000 899.500000 442.350000 ;
      RECT 807.500000 441.650000 849.500000 442.350000 ;
      RECT 757.500000 441.650000 799.500000 442.350000 ;
      RECT 707.500000 441.650000 733.500000 442.350000 ;
      RECT 657.500000 441.650000 699.500000 442.350000 ;
      RECT 607.500000 441.650000 649.500000 442.350000 ;
      RECT 557.500000 441.650000 599.500000 442.350000 ;
      RECT 507.500000 441.650000 549.500000 442.350000 ;
      RECT 457.500000 441.650000 499.500000 442.350000 ;
      RECT 407.500000 441.650000 449.500000 442.350000 ;
      RECT 357.500000 441.650000 399.500000 442.350000 ;
      RECT 307.500000 441.650000 349.500000 442.350000 ;
      RECT 207.500000 441.650000 299.500000 442.350000 ;
      RECT 107.500000 441.650000 199.500000 442.350000 ;
      RECT 57.500000 441.650000 99.500000 442.350000 ;
      RECT 15.500000 441.650000 49.500000 442.350000 ;
      RECT 1183.500000 440.350000 1186.000000 443.650000 ;
      RECT 1166.500000 440.350000 1170.500000 441.650000 ;
      RECT 1157.500000 440.350000 1158.500000 441.650000 ;
      RECT 1116.500000 440.350000 1149.500000 441.650000 ;
      RECT 1107.500000 440.350000 1108.500000 441.650000 ;
      RECT 1066.500000 440.350000 1099.500000 441.650000 ;
      RECT 1057.500000 440.350000 1058.500000 441.650000 ;
      RECT 1016.500000 440.350000 1049.500000 441.650000 ;
      RECT 1007.500000 440.350000 1008.500000 441.650000 ;
      RECT 966.500000 440.350000 999.500000 441.650000 ;
      RECT 957.500000 440.350000 958.500000 441.650000 ;
      RECT 916.500000 440.350000 949.500000 441.650000 ;
      RECT 907.500000 440.350000 908.500000 441.650000 ;
      RECT 866.500000 440.350000 899.500000 441.650000 ;
      RECT 857.500000 440.350000 858.500000 441.650000 ;
      RECT 816.500000 440.350000 849.500000 441.650000 ;
      RECT 807.500000 440.350000 808.500000 441.650000 ;
      RECT 766.500000 440.350000 799.500000 441.650000 ;
      RECT 757.500000 440.350000 758.500000 441.650000 ;
      RECT 746.500000 440.350000 749.500000 443.650000 ;
      RECT 732.500000 440.350000 733.500000 441.650000 ;
      RECT 707.500000 440.350000 708.500000 441.650000 ;
      RECT 666.500000 440.350000 699.500000 441.650000 ;
      RECT 657.500000 440.350000 658.500000 441.650000 ;
      RECT 616.500000 440.350000 649.500000 441.650000 ;
      RECT 607.500000 440.350000 608.500000 441.650000 ;
      RECT 566.500000 440.350000 599.500000 441.650000 ;
      RECT 557.500000 440.350000 558.500000 441.650000 ;
      RECT 516.500000 440.350000 549.500000 441.650000 ;
      RECT 507.500000 440.350000 508.500000 441.650000 ;
      RECT 466.500000 440.350000 499.500000 441.650000 ;
      RECT 457.500000 440.350000 458.500000 441.650000 ;
      RECT 416.500000 440.350000 449.500000 441.650000 ;
      RECT 407.500000 440.350000 408.500000 441.650000 ;
      RECT 366.500000 440.350000 399.500000 441.650000 ;
      RECT 357.500000 440.350000 358.500000 441.650000 ;
      RECT 316.500000 440.350000 349.500000 441.650000 ;
      RECT 307.500000 440.350000 308.500000 441.650000 ;
      RECT 216.500000 440.350000 299.500000 441.650000 ;
      RECT 207.500000 440.350000 208.500000 441.650000 ;
      RECT 116.500000 440.350000 199.500000 441.650000 ;
      RECT 107.500000 440.350000 108.500000 441.650000 ;
      RECT 66.500000 440.350000 99.500000 441.650000 ;
      RECT 57.500000 440.350000 58.500000 441.650000 ;
      RECT 29.500000 440.350000 49.500000 441.650000 ;
      RECT 15.500000 440.350000 16.500000 441.650000 ;
      RECT 0.000000 440.350000 2.500000 443.650000 ;
      RECT 1166.500000 439.650000 1186.000000 440.350000 ;
      RECT 1116.500000 439.650000 1158.500000 440.350000 ;
      RECT 1066.500000 439.650000 1108.500000 440.350000 ;
      RECT 1016.500000 439.650000 1058.500000 440.350000 ;
      RECT 966.500000 439.650000 1008.500000 440.350000 ;
      RECT 916.500000 439.650000 958.500000 440.350000 ;
      RECT 866.500000 439.650000 908.500000 440.350000 ;
      RECT 816.500000 439.650000 858.500000 440.350000 ;
      RECT 766.500000 439.650000 808.500000 440.350000 ;
      RECT 732.500000 439.650000 758.500000 440.350000 ;
      RECT 666.500000 439.650000 708.500000 440.350000 ;
      RECT 616.500000 439.650000 658.500000 440.350000 ;
      RECT 566.500000 439.650000 608.500000 440.350000 ;
      RECT 516.500000 439.650000 558.500000 440.350000 ;
      RECT 466.500000 439.650000 508.500000 440.350000 ;
      RECT 416.500000 439.650000 458.500000 440.350000 ;
      RECT 366.500000 439.650000 408.500000 440.350000 ;
      RECT 316.500000 439.650000 358.500000 440.350000 ;
      RECT 216.500000 439.650000 308.500000 440.350000 ;
      RECT 116.500000 439.650000 208.500000 440.350000 ;
      RECT 66.500000 439.650000 108.500000 440.350000 ;
      RECT 29.500000 439.650000 58.500000 440.350000 ;
      RECT 0.000000 439.650000 16.500000 440.350000 ;
      RECT 1166.500000 438.350000 1170.500000 439.650000 ;
      RECT 1157.500000 438.350000 1158.500000 439.650000 ;
      RECT 1116.500000 438.350000 1149.500000 439.650000 ;
      RECT 1107.500000 438.350000 1108.500000 439.650000 ;
      RECT 1066.500000 438.350000 1099.500000 439.650000 ;
      RECT 1057.500000 438.350000 1058.500000 439.650000 ;
      RECT 1016.500000 438.350000 1049.500000 439.650000 ;
      RECT 1007.500000 438.350000 1008.500000 439.650000 ;
      RECT 966.500000 438.350000 999.500000 439.650000 ;
      RECT 957.500000 438.350000 958.500000 439.650000 ;
      RECT 916.500000 438.350000 949.500000 439.650000 ;
      RECT 907.500000 438.350000 908.500000 439.650000 ;
      RECT 866.500000 438.350000 899.500000 439.650000 ;
      RECT 857.500000 438.350000 858.500000 439.650000 ;
      RECT 816.500000 438.350000 849.500000 439.650000 ;
      RECT 807.500000 438.350000 808.500000 439.650000 ;
      RECT 766.500000 438.350000 799.500000 439.650000 ;
      RECT 757.500000 438.350000 758.500000 439.650000 ;
      RECT 732.500000 438.350000 733.500000 439.650000 ;
      RECT 716.500000 438.350000 719.500000 441.650000 ;
      RECT 707.500000 438.350000 708.500000 439.650000 ;
      RECT 666.500000 438.350000 699.500000 439.650000 ;
      RECT 657.500000 438.350000 658.500000 439.650000 ;
      RECT 616.500000 438.350000 649.500000 439.650000 ;
      RECT 607.500000 438.350000 608.500000 439.650000 ;
      RECT 566.500000 438.350000 599.500000 439.650000 ;
      RECT 557.500000 438.350000 558.500000 439.650000 ;
      RECT 516.500000 438.350000 549.500000 439.650000 ;
      RECT 507.500000 438.350000 508.500000 439.650000 ;
      RECT 466.500000 438.350000 499.500000 439.650000 ;
      RECT 457.500000 438.350000 458.500000 439.650000 ;
      RECT 416.500000 438.350000 449.500000 439.650000 ;
      RECT 407.500000 438.350000 408.500000 439.650000 ;
      RECT 366.500000 438.350000 399.500000 439.650000 ;
      RECT 357.500000 438.350000 358.500000 439.650000 ;
      RECT 316.500000 438.350000 349.500000 439.650000 ;
      RECT 307.500000 438.350000 308.500000 439.650000 ;
      RECT 216.500000 438.350000 299.500000 439.650000 ;
      RECT 207.500000 438.350000 208.500000 439.650000 ;
      RECT 116.500000 438.350000 199.500000 439.650000 ;
      RECT 107.500000 438.350000 108.500000 439.650000 ;
      RECT 66.500000 438.350000 99.500000 439.650000 ;
      RECT 57.500000 438.350000 58.500000 439.650000 ;
      RECT 29.500000 438.350000 49.500000 439.650000 ;
      RECT 15.500000 438.350000 16.500000 439.650000 ;
      RECT 1157.500000 437.650000 1170.500000 438.350000 ;
      RECT 1107.500000 437.650000 1149.500000 438.350000 ;
      RECT 1057.500000 437.650000 1099.500000 438.350000 ;
      RECT 1007.500000 437.650000 1049.500000 438.350000 ;
      RECT 957.500000 437.650000 999.500000 438.350000 ;
      RECT 907.500000 437.650000 949.500000 438.350000 ;
      RECT 857.500000 437.650000 899.500000 438.350000 ;
      RECT 807.500000 437.650000 849.500000 438.350000 ;
      RECT 757.500000 437.650000 799.500000 438.350000 ;
      RECT 707.500000 437.650000 733.500000 438.350000 ;
      RECT 657.500000 437.650000 699.500000 438.350000 ;
      RECT 607.500000 437.650000 649.500000 438.350000 ;
      RECT 557.500000 437.650000 599.500000 438.350000 ;
      RECT 507.500000 437.650000 549.500000 438.350000 ;
      RECT 457.500000 437.650000 499.500000 438.350000 ;
      RECT 407.500000 437.650000 449.500000 438.350000 ;
      RECT 357.500000 437.650000 399.500000 438.350000 ;
      RECT 307.500000 437.650000 349.500000 438.350000 ;
      RECT 207.500000 437.650000 299.500000 438.350000 ;
      RECT 107.500000 437.650000 199.500000 438.350000 ;
      RECT 57.500000 437.650000 99.500000 438.350000 ;
      RECT 15.500000 437.650000 49.500000 438.350000 ;
      RECT 1183.500000 436.350000 1186.000000 439.650000 ;
      RECT 1166.500000 436.350000 1170.500000 437.650000 ;
      RECT 1157.500000 436.350000 1158.500000 437.650000 ;
      RECT 1116.500000 436.350000 1149.500000 437.650000 ;
      RECT 1107.500000 436.350000 1108.500000 437.650000 ;
      RECT 1066.500000 436.350000 1099.500000 437.650000 ;
      RECT 1057.500000 436.350000 1058.500000 437.650000 ;
      RECT 1016.500000 436.350000 1049.500000 437.650000 ;
      RECT 1007.500000 436.350000 1008.500000 437.650000 ;
      RECT 966.500000 436.350000 999.500000 437.650000 ;
      RECT 957.500000 436.350000 958.500000 437.650000 ;
      RECT 916.500000 436.350000 949.500000 437.650000 ;
      RECT 907.500000 436.350000 908.500000 437.650000 ;
      RECT 866.500000 436.350000 899.500000 437.650000 ;
      RECT 857.500000 436.350000 858.500000 437.650000 ;
      RECT 816.500000 436.350000 849.500000 437.650000 ;
      RECT 807.500000 436.350000 808.500000 437.650000 ;
      RECT 766.500000 436.350000 799.500000 437.650000 ;
      RECT 757.500000 436.350000 758.500000 437.650000 ;
      RECT 746.500000 436.350000 749.500000 439.650000 ;
      RECT 732.500000 436.350000 733.500000 437.650000 ;
      RECT 707.500000 436.350000 708.500000 437.650000 ;
      RECT 666.500000 436.350000 699.500000 437.650000 ;
      RECT 657.500000 436.350000 658.500000 437.650000 ;
      RECT 616.500000 436.350000 649.500000 437.650000 ;
      RECT 607.500000 436.350000 608.500000 437.650000 ;
      RECT 566.500000 436.350000 599.500000 437.650000 ;
      RECT 557.500000 436.350000 558.500000 437.650000 ;
      RECT 516.500000 436.350000 549.500000 437.650000 ;
      RECT 507.500000 436.350000 508.500000 437.650000 ;
      RECT 466.500000 436.350000 499.500000 437.650000 ;
      RECT 457.500000 436.350000 458.500000 437.650000 ;
      RECT 416.500000 436.350000 449.500000 437.650000 ;
      RECT 407.500000 436.350000 408.500000 437.650000 ;
      RECT 366.500000 436.350000 399.500000 437.650000 ;
      RECT 357.500000 436.350000 358.500000 437.650000 ;
      RECT 316.500000 436.350000 349.500000 437.650000 ;
      RECT 307.500000 436.350000 308.500000 437.650000 ;
      RECT 216.500000 436.350000 299.500000 437.650000 ;
      RECT 207.500000 436.350000 208.500000 437.650000 ;
      RECT 116.500000 436.350000 199.500000 437.650000 ;
      RECT 107.500000 436.350000 108.500000 437.650000 ;
      RECT 66.500000 436.350000 99.500000 437.650000 ;
      RECT 57.500000 436.350000 58.500000 437.650000 ;
      RECT 29.500000 436.350000 49.500000 437.650000 ;
      RECT 15.500000 436.350000 16.500000 437.650000 ;
      RECT 0.000000 436.350000 2.500000 439.650000 ;
      RECT 1166.500000 435.650000 1186.000000 436.350000 ;
      RECT 1116.500000 435.650000 1158.500000 436.350000 ;
      RECT 1066.500000 435.650000 1108.500000 436.350000 ;
      RECT 1016.500000 435.650000 1058.500000 436.350000 ;
      RECT 966.500000 435.650000 1008.500000 436.350000 ;
      RECT 916.500000 435.650000 958.500000 436.350000 ;
      RECT 866.500000 435.650000 908.500000 436.350000 ;
      RECT 816.500000 435.650000 858.500000 436.350000 ;
      RECT 766.500000 435.650000 808.500000 436.350000 ;
      RECT 732.500000 435.650000 758.500000 436.350000 ;
      RECT 666.500000 435.650000 708.500000 436.350000 ;
      RECT 616.500000 435.650000 658.500000 436.350000 ;
      RECT 566.500000 435.650000 608.500000 436.350000 ;
      RECT 516.500000 435.650000 558.500000 436.350000 ;
      RECT 466.500000 435.650000 508.500000 436.350000 ;
      RECT 416.500000 435.650000 458.500000 436.350000 ;
      RECT 366.500000 435.650000 408.500000 436.350000 ;
      RECT 316.500000 435.650000 358.500000 436.350000 ;
      RECT 216.500000 435.650000 308.500000 436.350000 ;
      RECT 116.500000 435.650000 208.500000 436.350000 ;
      RECT 66.500000 435.650000 108.500000 436.350000 ;
      RECT 29.500000 435.650000 58.500000 436.350000 ;
      RECT 0.000000 435.650000 16.500000 436.350000 ;
      RECT 1166.500000 434.350000 1170.500000 435.650000 ;
      RECT 1157.500000 434.350000 1158.500000 435.650000 ;
      RECT 1116.500000 434.350000 1149.500000 435.650000 ;
      RECT 1107.500000 434.350000 1108.500000 435.650000 ;
      RECT 1066.500000 434.350000 1099.500000 435.650000 ;
      RECT 1057.500000 434.350000 1058.500000 435.650000 ;
      RECT 1016.500000 434.350000 1049.500000 435.650000 ;
      RECT 1007.500000 434.350000 1008.500000 435.650000 ;
      RECT 966.500000 434.350000 999.500000 435.650000 ;
      RECT 957.500000 434.350000 958.500000 435.650000 ;
      RECT 916.500000 434.350000 949.500000 435.650000 ;
      RECT 907.500000 434.350000 908.500000 435.650000 ;
      RECT 866.500000 434.350000 899.500000 435.650000 ;
      RECT 857.500000 434.350000 858.500000 435.650000 ;
      RECT 816.500000 434.350000 849.500000 435.650000 ;
      RECT 807.500000 434.350000 808.500000 435.650000 ;
      RECT 766.500000 434.350000 799.500000 435.650000 ;
      RECT 757.500000 434.350000 758.500000 435.650000 ;
      RECT 732.500000 434.350000 733.500000 435.650000 ;
      RECT 716.500000 434.350000 719.500000 437.650000 ;
      RECT 707.500000 434.350000 708.500000 435.650000 ;
      RECT 666.500000 434.350000 699.500000 435.650000 ;
      RECT 657.500000 434.350000 658.500000 435.650000 ;
      RECT 616.500000 434.350000 649.500000 435.650000 ;
      RECT 607.500000 434.350000 608.500000 435.650000 ;
      RECT 566.500000 434.350000 599.500000 435.650000 ;
      RECT 557.500000 434.350000 558.500000 435.650000 ;
      RECT 516.500000 434.350000 549.500000 435.650000 ;
      RECT 507.500000 434.350000 508.500000 435.650000 ;
      RECT 466.500000 434.350000 499.500000 435.650000 ;
      RECT 457.500000 434.350000 458.500000 435.650000 ;
      RECT 416.500000 434.350000 449.500000 435.650000 ;
      RECT 407.500000 434.350000 408.500000 435.650000 ;
      RECT 366.500000 434.350000 399.500000 435.650000 ;
      RECT 357.500000 434.350000 358.500000 435.650000 ;
      RECT 316.500000 434.350000 349.500000 435.650000 ;
      RECT 307.500000 434.350000 308.500000 435.650000 ;
      RECT 216.500000 434.350000 299.500000 435.650000 ;
      RECT 207.500000 434.350000 208.500000 435.650000 ;
      RECT 116.500000 434.350000 199.500000 435.650000 ;
      RECT 107.500000 434.350000 108.500000 435.650000 ;
      RECT 66.500000 434.350000 99.500000 435.650000 ;
      RECT 57.500000 434.350000 58.500000 435.650000 ;
      RECT 29.500000 434.350000 49.500000 435.650000 ;
      RECT 15.500000 434.350000 16.500000 435.650000 ;
      RECT 1157.500000 433.650000 1170.500000 434.350000 ;
      RECT 1107.500000 433.650000 1149.500000 434.350000 ;
      RECT 1057.500000 433.650000 1099.500000 434.350000 ;
      RECT 1007.500000 433.650000 1049.500000 434.350000 ;
      RECT 957.500000 433.650000 999.500000 434.350000 ;
      RECT 907.500000 433.650000 949.500000 434.350000 ;
      RECT 857.500000 433.650000 899.500000 434.350000 ;
      RECT 807.500000 433.650000 849.500000 434.350000 ;
      RECT 757.500000 433.650000 799.500000 434.350000 ;
      RECT 707.500000 433.650000 733.500000 434.350000 ;
      RECT 657.500000 433.650000 699.500000 434.350000 ;
      RECT 607.500000 433.650000 649.500000 434.350000 ;
      RECT 557.500000 433.650000 599.500000 434.350000 ;
      RECT 507.500000 433.650000 549.500000 434.350000 ;
      RECT 457.500000 433.650000 499.500000 434.350000 ;
      RECT 407.500000 433.650000 449.500000 434.350000 ;
      RECT 357.500000 433.650000 399.500000 434.350000 ;
      RECT 307.500000 433.650000 349.500000 434.350000 ;
      RECT 207.500000 433.650000 299.500000 434.350000 ;
      RECT 107.500000 433.650000 199.500000 434.350000 ;
      RECT 57.500000 433.650000 99.500000 434.350000 ;
      RECT 15.500000 433.650000 49.500000 434.350000 ;
      RECT 1183.500000 432.350000 1186.000000 435.650000 ;
      RECT 1166.500000 432.350000 1170.500000 433.650000 ;
      RECT 1157.500000 432.350000 1158.500000 433.650000 ;
      RECT 1116.500000 432.350000 1149.500000 433.650000 ;
      RECT 1107.500000 432.350000 1108.500000 433.650000 ;
      RECT 1066.500000 432.350000 1099.500000 433.650000 ;
      RECT 1057.500000 432.350000 1058.500000 433.650000 ;
      RECT 1016.500000 432.350000 1049.500000 433.650000 ;
      RECT 1007.500000 432.350000 1008.500000 433.650000 ;
      RECT 966.500000 432.350000 999.500000 433.650000 ;
      RECT 957.500000 432.350000 958.500000 433.650000 ;
      RECT 916.500000 432.350000 949.500000 433.650000 ;
      RECT 907.500000 432.350000 908.500000 433.650000 ;
      RECT 866.500000 432.350000 899.500000 433.650000 ;
      RECT 857.500000 432.350000 858.500000 433.650000 ;
      RECT 816.500000 432.350000 849.500000 433.650000 ;
      RECT 807.500000 432.350000 808.500000 433.650000 ;
      RECT 766.500000 432.350000 799.500000 433.650000 ;
      RECT 757.500000 432.350000 758.500000 433.650000 ;
      RECT 746.500000 432.350000 749.500000 435.650000 ;
      RECT 732.500000 432.350000 733.500000 433.650000 ;
      RECT 707.500000 432.350000 708.500000 433.650000 ;
      RECT 666.500000 432.350000 699.500000 433.650000 ;
      RECT 657.500000 432.350000 658.500000 433.650000 ;
      RECT 616.500000 432.350000 649.500000 433.650000 ;
      RECT 607.500000 432.350000 608.500000 433.650000 ;
      RECT 566.500000 432.350000 599.500000 433.650000 ;
      RECT 557.500000 432.350000 558.500000 433.650000 ;
      RECT 516.500000 432.350000 549.500000 433.650000 ;
      RECT 507.500000 432.350000 508.500000 433.650000 ;
      RECT 466.500000 432.350000 499.500000 433.650000 ;
      RECT 457.500000 432.350000 458.500000 433.650000 ;
      RECT 416.500000 432.350000 449.500000 433.650000 ;
      RECT 407.500000 432.350000 408.500000 433.650000 ;
      RECT 366.500000 432.350000 399.500000 433.650000 ;
      RECT 357.500000 432.350000 358.500000 433.650000 ;
      RECT 316.500000 432.350000 349.500000 433.650000 ;
      RECT 307.500000 432.350000 308.500000 433.650000 ;
      RECT 216.500000 432.350000 299.500000 433.650000 ;
      RECT 207.500000 432.350000 208.500000 433.650000 ;
      RECT 116.500000 432.350000 199.500000 433.650000 ;
      RECT 107.500000 432.350000 108.500000 433.650000 ;
      RECT 66.500000 432.350000 99.500000 433.650000 ;
      RECT 57.500000 432.350000 58.500000 433.650000 ;
      RECT 29.500000 432.350000 49.500000 433.650000 ;
      RECT 15.500000 432.350000 16.500000 433.650000 ;
      RECT 0.000000 432.350000 2.500000 435.650000 ;
      RECT 1166.500000 431.650000 1186.000000 432.350000 ;
      RECT 1116.500000 431.650000 1158.500000 432.350000 ;
      RECT 1066.500000 431.650000 1108.500000 432.350000 ;
      RECT 1016.500000 431.650000 1058.500000 432.350000 ;
      RECT 966.500000 431.650000 1008.500000 432.350000 ;
      RECT 916.500000 431.650000 958.500000 432.350000 ;
      RECT 866.500000 431.650000 908.500000 432.350000 ;
      RECT 816.500000 431.650000 858.500000 432.350000 ;
      RECT 766.500000 431.650000 808.500000 432.350000 ;
      RECT 732.500000 431.650000 758.500000 432.350000 ;
      RECT 666.500000 431.650000 708.500000 432.350000 ;
      RECT 616.500000 431.650000 658.500000 432.350000 ;
      RECT 566.500000 431.650000 608.500000 432.350000 ;
      RECT 516.500000 431.650000 558.500000 432.350000 ;
      RECT 466.500000 431.650000 508.500000 432.350000 ;
      RECT 416.500000 431.650000 458.500000 432.350000 ;
      RECT 366.500000 431.650000 408.500000 432.350000 ;
      RECT 316.500000 431.650000 358.500000 432.350000 ;
      RECT 216.500000 431.650000 308.500000 432.350000 ;
      RECT 116.500000 431.650000 208.500000 432.350000 ;
      RECT 66.500000 431.650000 108.500000 432.350000 ;
      RECT 29.500000 431.650000 58.500000 432.350000 ;
      RECT 0.000000 431.650000 16.500000 432.350000 ;
      RECT 1166.500000 430.350000 1170.500000 431.650000 ;
      RECT 1157.500000 430.350000 1158.500000 431.650000 ;
      RECT 1116.500000 430.350000 1149.500000 431.650000 ;
      RECT 1107.500000 430.350000 1108.500000 431.650000 ;
      RECT 1066.500000 430.350000 1099.500000 431.650000 ;
      RECT 1057.500000 430.350000 1058.500000 431.650000 ;
      RECT 1016.500000 430.350000 1049.500000 431.650000 ;
      RECT 1007.500000 430.350000 1008.500000 431.650000 ;
      RECT 966.500000 430.350000 999.500000 431.650000 ;
      RECT 957.500000 430.350000 958.500000 431.650000 ;
      RECT 916.500000 430.350000 949.500000 431.650000 ;
      RECT 907.500000 430.350000 908.500000 431.650000 ;
      RECT 866.500000 430.350000 899.500000 431.650000 ;
      RECT 857.500000 430.350000 858.500000 431.650000 ;
      RECT 816.500000 430.350000 849.500000 431.650000 ;
      RECT 807.500000 430.350000 808.500000 431.650000 ;
      RECT 766.500000 430.350000 799.500000 431.650000 ;
      RECT 757.500000 430.350000 758.500000 431.650000 ;
      RECT 732.500000 430.350000 749.500000 431.650000 ;
      RECT 716.500000 430.350000 719.500000 433.650000 ;
      RECT 707.500000 430.350000 708.500000 431.650000 ;
      RECT 666.500000 430.350000 699.500000 431.650000 ;
      RECT 657.500000 430.350000 658.500000 431.650000 ;
      RECT 616.500000 430.350000 649.500000 431.650000 ;
      RECT 607.500000 430.350000 608.500000 431.650000 ;
      RECT 566.500000 430.350000 599.500000 431.650000 ;
      RECT 557.500000 430.350000 558.500000 431.650000 ;
      RECT 516.500000 430.350000 549.500000 431.650000 ;
      RECT 507.500000 430.350000 508.500000 431.650000 ;
      RECT 466.500000 430.350000 499.500000 431.650000 ;
      RECT 457.500000 430.350000 458.500000 431.650000 ;
      RECT 416.500000 430.350000 449.500000 431.650000 ;
      RECT 407.500000 430.350000 408.500000 431.650000 ;
      RECT 366.500000 430.350000 399.500000 431.650000 ;
      RECT 357.500000 430.350000 358.500000 431.650000 ;
      RECT 316.500000 430.350000 349.500000 431.650000 ;
      RECT 307.500000 430.350000 308.500000 431.650000 ;
      RECT 216.500000 430.350000 299.500000 431.650000 ;
      RECT 207.500000 430.350000 208.500000 431.650000 ;
      RECT 116.500000 430.350000 199.500000 431.650000 ;
      RECT 107.500000 430.350000 108.500000 431.650000 ;
      RECT 66.500000 430.350000 99.500000 431.650000 ;
      RECT 57.500000 430.350000 58.500000 431.650000 ;
      RECT 29.500000 430.350000 49.500000 431.650000 ;
      RECT 15.500000 430.350000 16.500000 431.650000 ;
      RECT 1157.500000 429.650000 1170.500000 430.350000 ;
      RECT 1107.500000 429.650000 1149.500000 430.350000 ;
      RECT 1057.500000 429.650000 1099.500000 430.350000 ;
      RECT 1007.500000 429.650000 1049.500000 430.350000 ;
      RECT 957.500000 429.650000 999.500000 430.350000 ;
      RECT 907.500000 429.650000 949.500000 430.350000 ;
      RECT 857.500000 429.650000 899.500000 430.350000 ;
      RECT 807.500000 429.650000 849.500000 430.350000 ;
      RECT 757.500000 429.650000 799.500000 430.350000 ;
      RECT 707.500000 429.650000 749.500000 430.350000 ;
      RECT 657.500000 429.650000 699.500000 430.350000 ;
      RECT 607.500000 429.650000 649.500000 430.350000 ;
      RECT 557.500000 429.650000 599.500000 430.350000 ;
      RECT 507.500000 429.650000 549.500000 430.350000 ;
      RECT 457.500000 429.650000 499.500000 430.350000 ;
      RECT 407.500000 429.650000 449.500000 430.350000 ;
      RECT 357.500000 429.650000 399.500000 430.350000 ;
      RECT 307.500000 429.650000 349.500000 430.350000 ;
      RECT 207.500000 429.650000 299.500000 430.350000 ;
      RECT 107.500000 429.650000 199.500000 430.350000 ;
      RECT 57.500000 429.650000 99.500000 430.350000 ;
      RECT 15.500000 429.650000 49.500000 430.350000 ;
      RECT 1183.500000 428.350000 1186.000000 431.650000 ;
      RECT 1169.500000 428.350000 1170.500000 429.650000 ;
      RECT 1116.500000 428.350000 1149.500000 429.650000 ;
      RECT 1107.500000 428.350000 1108.500000 429.650000 ;
      RECT 1066.500000 428.350000 1099.500000 429.650000 ;
      RECT 1057.500000 428.350000 1058.500000 429.650000 ;
      RECT 1016.500000 428.350000 1049.500000 429.650000 ;
      RECT 1007.500000 428.350000 1008.500000 429.650000 ;
      RECT 966.500000 428.350000 999.500000 429.650000 ;
      RECT 957.500000 428.350000 958.500000 429.650000 ;
      RECT 916.500000 428.350000 949.500000 429.650000 ;
      RECT 907.500000 428.350000 908.500000 429.650000 ;
      RECT 866.500000 428.350000 899.500000 429.650000 ;
      RECT 857.500000 428.350000 858.500000 429.650000 ;
      RECT 816.500000 428.350000 849.500000 429.650000 ;
      RECT 807.500000 428.350000 808.500000 429.650000 ;
      RECT 766.500000 428.350000 799.500000 429.650000 ;
      RECT 757.500000 428.350000 758.500000 429.650000 ;
      RECT 732.500000 428.350000 749.500000 429.650000 ;
      RECT 707.500000 428.350000 708.500000 429.650000 ;
      RECT 666.500000 428.350000 699.500000 429.650000 ;
      RECT 657.500000 428.350000 658.500000 429.650000 ;
      RECT 616.500000 428.350000 649.500000 429.650000 ;
      RECT 607.500000 428.350000 608.500000 429.650000 ;
      RECT 566.500000 428.350000 599.500000 429.650000 ;
      RECT 557.500000 428.350000 558.500000 429.650000 ;
      RECT 516.500000 428.350000 549.500000 429.650000 ;
      RECT 507.500000 428.350000 508.500000 429.650000 ;
      RECT 466.500000 428.350000 499.500000 429.650000 ;
      RECT 457.500000 428.350000 458.500000 429.650000 ;
      RECT 416.500000 428.350000 449.500000 429.650000 ;
      RECT 407.500000 428.350000 408.500000 429.650000 ;
      RECT 366.500000 428.350000 399.500000 429.650000 ;
      RECT 357.500000 428.350000 358.500000 429.650000 ;
      RECT 316.500000 428.350000 349.500000 429.650000 ;
      RECT 307.500000 428.350000 308.500000 429.650000 ;
      RECT 216.500000 428.350000 299.500000 429.650000 ;
      RECT 207.500000 428.350000 208.500000 429.650000 ;
      RECT 116.500000 428.350000 199.500000 429.650000 ;
      RECT 107.500000 428.350000 108.500000 429.650000 ;
      RECT 66.500000 428.350000 99.500000 429.650000 ;
      RECT 57.500000 428.350000 58.500000 429.650000 ;
      RECT 29.500000 428.350000 49.500000 429.650000 ;
      RECT 15.500000 428.350000 16.500000 429.650000 ;
      RECT 0.000000 428.350000 2.500000 431.650000 ;
      RECT 1169.500000 427.650000 1186.000000 428.350000 ;
      RECT 1116.500000 427.650000 1156.500000 428.350000 ;
      RECT 1066.500000 427.650000 1108.500000 428.350000 ;
      RECT 1016.500000 427.650000 1058.500000 428.350000 ;
      RECT 966.500000 427.650000 1008.500000 428.350000 ;
      RECT 916.500000 427.650000 958.500000 428.350000 ;
      RECT 866.500000 427.650000 908.500000 428.350000 ;
      RECT 816.500000 427.650000 858.500000 428.350000 ;
      RECT 766.500000 427.650000 808.500000 428.350000 ;
      RECT 732.500000 427.650000 758.500000 428.350000 ;
      RECT 666.500000 427.650000 708.500000 428.350000 ;
      RECT 616.500000 427.650000 658.500000 428.350000 ;
      RECT 566.500000 427.650000 608.500000 428.350000 ;
      RECT 516.500000 427.650000 558.500000 428.350000 ;
      RECT 466.500000 427.650000 508.500000 428.350000 ;
      RECT 416.500000 427.650000 458.500000 428.350000 ;
      RECT 366.500000 427.650000 408.500000 428.350000 ;
      RECT 316.500000 427.650000 358.500000 428.350000 ;
      RECT 216.500000 427.650000 308.500000 428.350000 ;
      RECT 116.500000 427.650000 208.500000 428.350000 ;
      RECT 66.500000 427.650000 108.500000 428.350000 ;
      RECT 29.500000 427.650000 58.500000 428.350000 ;
      RECT 0.000000 427.650000 16.500000 428.350000 ;
      RECT 1169.500000 426.350000 1170.500000 427.650000 ;
      RECT 1116.500000 426.350000 1149.500000 427.650000 ;
      RECT 1107.500000 426.350000 1108.500000 427.650000 ;
      RECT 1066.500000 426.350000 1099.500000 427.650000 ;
      RECT 1057.500000 426.350000 1058.500000 427.650000 ;
      RECT 1016.500000 426.350000 1049.500000 427.650000 ;
      RECT 1007.500000 426.350000 1008.500000 427.650000 ;
      RECT 966.500000 426.350000 999.500000 427.650000 ;
      RECT 957.500000 426.350000 958.500000 427.650000 ;
      RECT 916.500000 426.350000 949.500000 427.650000 ;
      RECT 907.500000 426.350000 908.500000 427.650000 ;
      RECT 866.500000 426.350000 899.500000 427.650000 ;
      RECT 857.500000 426.350000 858.500000 427.650000 ;
      RECT 816.500000 426.350000 849.500000 427.650000 ;
      RECT 807.500000 426.350000 808.500000 427.650000 ;
      RECT 766.500000 426.350000 799.500000 427.650000 ;
      RECT 757.500000 426.350000 758.500000 427.650000 ;
      RECT 732.500000 426.350000 749.500000 427.650000 ;
      RECT 716.500000 426.350000 719.500000 429.650000 ;
      RECT 707.500000 426.350000 708.500000 427.650000 ;
      RECT 666.500000 426.350000 699.500000 427.650000 ;
      RECT 657.500000 426.350000 658.500000 427.650000 ;
      RECT 616.500000 426.350000 649.500000 427.650000 ;
      RECT 607.500000 426.350000 608.500000 427.650000 ;
      RECT 566.500000 426.350000 599.500000 427.650000 ;
      RECT 557.500000 426.350000 558.500000 427.650000 ;
      RECT 516.500000 426.350000 549.500000 427.650000 ;
      RECT 507.500000 426.350000 508.500000 427.650000 ;
      RECT 466.500000 426.350000 499.500000 427.650000 ;
      RECT 457.500000 426.350000 458.500000 427.650000 ;
      RECT 416.500000 426.350000 449.500000 427.650000 ;
      RECT 407.500000 426.350000 408.500000 427.650000 ;
      RECT 366.500000 426.350000 399.500000 427.650000 ;
      RECT 357.500000 426.350000 358.500000 427.650000 ;
      RECT 316.500000 426.350000 349.500000 427.650000 ;
      RECT 307.500000 426.350000 308.500000 427.650000 ;
      RECT 216.500000 426.350000 299.500000 427.650000 ;
      RECT 207.500000 426.350000 208.500000 427.650000 ;
      RECT 116.500000 426.350000 199.500000 427.650000 ;
      RECT 107.500000 426.350000 108.500000 427.650000 ;
      RECT 66.500000 426.350000 99.500000 427.650000 ;
      RECT 57.500000 426.350000 58.500000 427.650000 ;
      RECT 29.500000 426.350000 49.500000 427.650000 ;
      RECT 15.500000 426.350000 16.500000 427.650000 ;
      RECT 1157.500000 425.650000 1170.500000 426.350000 ;
      RECT 1107.500000 425.650000 1149.500000 426.350000 ;
      RECT 1057.500000 425.650000 1099.500000 426.350000 ;
      RECT 1007.500000 425.650000 1049.500000 426.350000 ;
      RECT 957.500000 425.650000 999.500000 426.350000 ;
      RECT 907.500000 425.650000 949.500000 426.350000 ;
      RECT 857.500000 425.650000 899.500000 426.350000 ;
      RECT 807.500000 425.650000 849.500000 426.350000 ;
      RECT 757.500000 425.650000 799.500000 426.350000 ;
      RECT 707.500000 425.650000 749.500000 426.350000 ;
      RECT 657.500000 425.650000 699.500000 426.350000 ;
      RECT 607.500000 425.650000 649.500000 426.350000 ;
      RECT 557.500000 425.650000 599.500000 426.350000 ;
      RECT 507.500000 425.650000 549.500000 426.350000 ;
      RECT 457.500000 425.650000 499.500000 426.350000 ;
      RECT 407.500000 425.650000 449.500000 426.350000 ;
      RECT 357.500000 425.650000 399.500000 426.350000 ;
      RECT 307.500000 425.650000 349.500000 426.350000 ;
      RECT 207.500000 425.650000 299.500000 426.350000 ;
      RECT 107.500000 425.650000 199.500000 426.350000 ;
      RECT 57.500000 425.650000 99.500000 426.350000 ;
      RECT 15.500000 425.650000 49.500000 426.350000 ;
      RECT 1183.500000 424.350000 1186.000000 427.650000 ;
      RECT 1169.500000 424.350000 1170.500000 425.650000 ;
      RECT 1116.500000 424.350000 1149.500000 425.650000 ;
      RECT 1107.500000 424.350000 1108.500000 425.650000 ;
      RECT 1066.500000 424.350000 1099.500000 425.650000 ;
      RECT 1057.500000 424.350000 1058.500000 425.650000 ;
      RECT 1016.500000 424.350000 1049.500000 425.650000 ;
      RECT 1007.500000 424.350000 1008.500000 425.650000 ;
      RECT 966.500000 424.350000 999.500000 425.650000 ;
      RECT 957.500000 424.350000 958.500000 425.650000 ;
      RECT 916.500000 424.350000 949.500000 425.650000 ;
      RECT 907.500000 424.350000 908.500000 425.650000 ;
      RECT 866.500000 424.350000 899.500000 425.650000 ;
      RECT 857.500000 424.350000 858.500000 425.650000 ;
      RECT 816.500000 424.350000 849.500000 425.650000 ;
      RECT 807.500000 424.350000 808.500000 425.650000 ;
      RECT 766.500000 424.350000 799.500000 425.650000 ;
      RECT 757.500000 424.350000 758.500000 425.650000 ;
      RECT 732.500000 424.350000 749.500000 425.650000 ;
      RECT 707.500000 424.350000 708.500000 425.650000 ;
      RECT 666.500000 424.350000 699.500000 425.650000 ;
      RECT 657.500000 424.350000 658.500000 425.650000 ;
      RECT 616.500000 424.350000 649.500000 425.650000 ;
      RECT 607.500000 424.350000 608.500000 425.650000 ;
      RECT 566.500000 424.350000 599.500000 425.650000 ;
      RECT 557.500000 424.350000 558.500000 425.650000 ;
      RECT 516.500000 424.350000 549.500000 425.650000 ;
      RECT 507.500000 424.350000 508.500000 425.650000 ;
      RECT 466.500000 424.350000 499.500000 425.650000 ;
      RECT 457.500000 424.350000 458.500000 425.650000 ;
      RECT 416.500000 424.350000 449.500000 425.650000 ;
      RECT 407.500000 424.350000 408.500000 425.650000 ;
      RECT 366.500000 424.350000 399.500000 425.650000 ;
      RECT 357.500000 424.350000 358.500000 425.650000 ;
      RECT 316.500000 424.350000 349.500000 425.650000 ;
      RECT 307.500000 424.350000 308.500000 425.650000 ;
      RECT 216.500000 424.350000 299.500000 425.650000 ;
      RECT 207.500000 424.350000 208.500000 425.650000 ;
      RECT 116.500000 424.350000 199.500000 425.650000 ;
      RECT 107.500000 424.350000 108.500000 425.650000 ;
      RECT 66.500000 424.350000 99.500000 425.650000 ;
      RECT 57.500000 424.350000 58.500000 425.650000 ;
      RECT 29.500000 424.350000 49.500000 425.650000 ;
      RECT 15.500000 424.350000 16.500000 425.650000 ;
      RECT 0.000000 424.350000 2.500000 427.650000 ;
      RECT 1169.500000 423.650000 1186.000000 424.350000 ;
      RECT 1116.500000 423.650000 1156.500000 424.350000 ;
      RECT 1066.500000 423.650000 1108.500000 424.350000 ;
      RECT 1016.500000 423.650000 1058.500000 424.350000 ;
      RECT 966.500000 423.650000 1008.500000 424.350000 ;
      RECT 916.500000 423.650000 958.500000 424.350000 ;
      RECT 866.500000 423.650000 908.500000 424.350000 ;
      RECT 816.500000 423.650000 858.500000 424.350000 ;
      RECT 766.500000 423.650000 808.500000 424.350000 ;
      RECT 732.500000 423.650000 758.500000 424.350000 ;
      RECT 666.500000 423.650000 708.500000 424.350000 ;
      RECT 616.500000 423.650000 658.500000 424.350000 ;
      RECT 566.500000 423.650000 608.500000 424.350000 ;
      RECT 516.500000 423.650000 558.500000 424.350000 ;
      RECT 466.500000 423.650000 508.500000 424.350000 ;
      RECT 416.500000 423.650000 458.500000 424.350000 ;
      RECT 366.500000 423.650000 408.500000 424.350000 ;
      RECT 316.500000 423.650000 358.500000 424.350000 ;
      RECT 216.500000 423.650000 308.500000 424.350000 ;
      RECT 116.500000 423.650000 208.500000 424.350000 ;
      RECT 66.500000 423.650000 108.500000 424.350000 ;
      RECT 29.500000 423.650000 58.500000 424.350000 ;
      RECT 0.000000 423.650000 16.500000 424.350000 ;
      RECT 1169.500000 422.350000 1170.500000 423.650000 ;
      RECT 1116.500000 422.350000 1149.500000 423.650000 ;
      RECT 1107.500000 422.350000 1108.500000 423.650000 ;
      RECT 1066.500000 422.350000 1099.500000 423.650000 ;
      RECT 1057.500000 422.350000 1058.500000 423.650000 ;
      RECT 1016.500000 422.350000 1049.500000 423.650000 ;
      RECT 1007.500000 422.350000 1008.500000 423.650000 ;
      RECT 966.500000 422.350000 999.500000 423.650000 ;
      RECT 957.500000 422.350000 958.500000 423.650000 ;
      RECT 916.500000 422.350000 949.500000 423.650000 ;
      RECT 907.500000 422.350000 908.500000 423.650000 ;
      RECT 866.500000 422.350000 899.500000 423.650000 ;
      RECT 857.500000 422.350000 858.500000 423.650000 ;
      RECT 816.500000 422.350000 849.500000 423.650000 ;
      RECT 807.500000 422.350000 808.500000 423.650000 ;
      RECT 766.500000 422.350000 799.500000 423.650000 ;
      RECT 757.500000 422.350000 758.500000 423.650000 ;
      RECT 732.500000 422.350000 749.500000 423.650000 ;
      RECT 716.500000 422.350000 719.500000 425.650000 ;
      RECT 707.500000 422.350000 708.500000 423.650000 ;
      RECT 666.500000 422.350000 699.500000 423.650000 ;
      RECT 657.500000 422.350000 658.500000 423.650000 ;
      RECT 616.500000 422.350000 649.500000 423.650000 ;
      RECT 607.500000 422.350000 608.500000 423.650000 ;
      RECT 566.500000 422.350000 599.500000 423.650000 ;
      RECT 557.500000 422.350000 558.500000 423.650000 ;
      RECT 516.500000 422.350000 549.500000 423.650000 ;
      RECT 507.500000 422.350000 508.500000 423.650000 ;
      RECT 466.500000 422.350000 499.500000 423.650000 ;
      RECT 457.500000 422.350000 458.500000 423.650000 ;
      RECT 416.500000 422.350000 449.500000 423.650000 ;
      RECT 407.500000 422.350000 408.500000 423.650000 ;
      RECT 366.500000 422.350000 399.500000 423.650000 ;
      RECT 357.500000 422.350000 358.500000 423.650000 ;
      RECT 316.500000 422.350000 349.500000 423.650000 ;
      RECT 307.500000 422.350000 308.500000 423.650000 ;
      RECT 216.500000 422.350000 299.500000 423.650000 ;
      RECT 207.500000 422.350000 208.500000 423.650000 ;
      RECT 116.500000 422.350000 199.500000 423.650000 ;
      RECT 107.500000 422.350000 108.500000 423.650000 ;
      RECT 66.500000 422.350000 99.500000 423.650000 ;
      RECT 57.500000 422.350000 58.500000 423.650000 ;
      RECT 29.500000 422.350000 49.500000 423.650000 ;
      RECT 15.500000 422.350000 16.500000 423.650000 ;
      RECT 1157.500000 421.650000 1170.500000 422.350000 ;
      RECT 1107.500000 421.650000 1149.500000 422.350000 ;
      RECT 1057.500000 421.650000 1099.500000 422.350000 ;
      RECT 1007.500000 421.650000 1049.500000 422.350000 ;
      RECT 957.500000 421.650000 999.500000 422.350000 ;
      RECT 907.500000 421.650000 949.500000 422.350000 ;
      RECT 857.500000 421.650000 899.500000 422.350000 ;
      RECT 807.500000 421.650000 849.500000 422.350000 ;
      RECT 757.500000 421.650000 799.500000 422.350000 ;
      RECT 707.500000 421.650000 749.500000 422.350000 ;
      RECT 657.500000 421.650000 699.500000 422.350000 ;
      RECT 607.500000 421.650000 649.500000 422.350000 ;
      RECT 557.500000 421.650000 599.500000 422.350000 ;
      RECT 507.500000 421.650000 549.500000 422.350000 ;
      RECT 457.500000 421.650000 499.500000 422.350000 ;
      RECT 407.500000 421.650000 449.500000 422.350000 ;
      RECT 357.500000 421.650000 399.500000 422.350000 ;
      RECT 307.500000 421.650000 349.500000 422.350000 ;
      RECT 207.500000 421.650000 299.500000 422.350000 ;
      RECT 107.500000 421.650000 199.500000 422.350000 ;
      RECT 57.500000 421.650000 99.500000 422.350000 ;
      RECT 15.500000 421.650000 49.500000 422.350000 ;
      RECT 1183.500000 420.350000 1186.000000 423.650000 ;
      RECT 1169.500000 420.350000 1170.500000 421.650000 ;
      RECT 1116.500000 420.350000 1149.500000 421.650000 ;
      RECT 1107.500000 420.350000 1108.500000 421.650000 ;
      RECT 1066.500000 420.350000 1099.500000 421.650000 ;
      RECT 1057.500000 420.350000 1058.500000 421.650000 ;
      RECT 1016.500000 420.350000 1049.500000 421.650000 ;
      RECT 1007.500000 420.350000 1008.500000 421.650000 ;
      RECT 966.500000 420.350000 999.500000 421.650000 ;
      RECT 957.500000 420.350000 958.500000 421.650000 ;
      RECT 916.500000 420.350000 949.500000 421.650000 ;
      RECT 907.500000 420.350000 908.500000 421.650000 ;
      RECT 866.500000 420.350000 899.500000 421.650000 ;
      RECT 857.500000 420.350000 858.500000 421.650000 ;
      RECT 816.500000 420.350000 849.500000 421.650000 ;
      RECT 807.500000 420.350000 808.500000 421.650000 ;
      RECT 766.500000 420.350000 799.500000 421.650000 ;
      RECT 757.500000 420.350000 758.500000 421.650000 ;
      RECT 732.500000 420.350000 749.500000 421.650000 ;
      RECT 707.500000 420.350000 708.500000 421.650000 ;
      RECT 666.500000 420.350000 699.500000 421.650000 ;
      RECT 657.500000 420.350000 658.500000 421.650000 ;
      RECT 616.500000 420.350000 649.500000 421.650000 ;
      RECT 607.500000 420.350000 608.500000 421.650000 ;
      RECT 566.500000 420.350000 599.500000 421.650000 ;
      RECT 557.500000 420.350000 558.500000 421.650000 ;
      RECT 516.500000 420.350000 549.500000 421.650000 ;
      RECT 507.500000 420.350000 508.500000 421.650000 ;
      RECT 466.500000 420.350000 499.500000 421.650000 ;
      RECT 457.500000 420.350000 458.500000 421.650000 ;
      RECT 416.500000 420.350000 449.500000 421.650000 ;
      RECT 407.500000 420.350000 408.500000 421.650000 ;
      RECT 366.500000 420.350000 399.500000 421.650000 ;
      RECT 357.500000 420.350000 358.500000 421.650000 ;
      RECT 316.500000 420.350000 349.500000 421.650000 ;
      RECT 307.500000 420.350000 308.500000 421.650000 ;
      RECT 216.500000 420.350000 299.500000 421.650000 ;
      RECT 207.500000 420.350000 208.500000 421.650000 ;
      RECT 116.500000 420.350000 199.500000 421.650000 ;
      RECT 107.500000 420.350000 108.500000 421.650000 ;
      RECT 66.500000 420.350000 99.500000 421.650000 ;
      RECT 57.500000 420.350000 58.500000 421.650000 ;
      RECT 29.500000 420.350000 49.500000 421.650000 ;
      RECT 15.500000 420.350000 16.500000 421.650000 ;
      RECT 0.000000 420.350000 2.500000 423.650000 ;
      RECT 1169.500000 419.650000 1186.000000 420.350000 ;
      RECT 1116.500000 419.650000 1156.500000 420.350000 ;
      RECT 1066.500000 419.650000 1108.500000 420.350000 ;
      RECT 1016.500000 419.650000 1058.500000 420.350000 ;
      RECT 966.500000 419.650000 1008.500000 420.350000 ;
      RECT 916.500000 419.650000 958.500000 420.350000 ;
      RECT 866.500000 419.650000 908.500000 420.350000 ;
      RECT 816.500000 419.650000 858.500000 420.350000 ;
      RECT 766.500000 419.650000 808.500000 420.350000 ;
      RECT 732.500000 419.650000 758.500000 420.350000 ;
      RECT 666.500000 419.650000 708.500000 420.350000 ;
      RECT 616.500000 419.650000 658.500000 420.350000 ;
      RECT 566.500000 419.650000 608.500000 420.350000 ;
      RECT 516.500000 419.650000 558.500000 420.350000 ;
      RECT 466.500000 419.650000 508.500000 420.350000 ;
      RECT 366.500000 419.650000 408.500000 420.350000 ;
      RECT 316.500000 419.650000 358.500000 420.350000 ;
      RECT 216.500000 419.650000 308.500000 420.350000 ;
      RECT 116.500000 419.650000 208.500000 420.350000 ;
      RECT 66.500000 419.650000 108.500000 420.350000 ;
      RECT 29.500000 419.650000 58.500000 420.350000 ;
      RECT 0.000000 419.650000 16.500000 420.350000 ;
      RECT 1169.500000 418.350000 1170.500000 419.650000 ;
      RECT 1116.500000 418.350000 1149.500000 419.650000 ;
      RECT 1107.500000 418.350000 1108.500000 419.650000 ;
      RECT 1066.500000 418.350000 1099.500000 419.650000 ;
      RECT 1057.500000 418.350000 1058.500000 419.650000 ;
      RECT 1016.500000 418.350000 1049.500000 419.650000 ;
      RECT 1007.500000 418.350000 1008.500000 419.650000 ;
      RECT 966.500000 418.350000 999.500000 419.650000 ;
      RECT 957.500000 418.350000 958.500000 419.650000 ;
      RECT 916.500000 418.350000 949.500000 419.650000 ;
      RECT 907.500000 418.350000 908.500000 419.650000 ;
      RECT 866.500000 418.350000 899.500000 419.650000 ;
      RECT 857.500000 418.350000 858.500000 419.650000 ;
      RECT 816.500000 418.350000 849.500000 419.650000 ;
      RECT 807.500000 418.350000 808.500000 419.650000 ;
      RECT 766.500000 418.350000 799.500000 419.650000 ;
      RECT 757.500000 418.350000 758.500000 419.650000 ;
      RECT 732.500000 418.350000 749.500000 419.650000 ;
      RECT 716.500000 418.350000 719.500000 421.650000 ;
      RECT 707.500000 418.350000 708.500000 419.650000 ;
      RECT 666.500000 418.350000 699.500000 419.650000 ;
      RECT 657.500000 418.350000 658.500000 419.650000 ;
      RECT 616.500000 418.350000 649.500000 419.650000 ;
      RECT 607.500000 418.350000 608.500000 419.650000 ;
      RECT 566.500000 418.350000 599.500000 419.650000 ;
      RECT 557.500000 418.350000 558.500000 419.650000 ;
      RECT 516.500000 418.350000 549.500000 419.650000 ;
      RECT 507.500000 418.350000 508.500000 419.650000 ;
      RECT 466.500000 418.350000 499.500000 419.650000 ;
      RECT 416.500000 418.350000 458.500000 420.350000 ;
      RECT 407.500000 418.350000 408.500000 419.650000 ;
      RECT 366.500000 418.350000 399.500000 419.650000 ;
      RECT 357.500000 418.350000 358.500000 419.650000 ;
      RECT 316.500000 418.350000 349.500000 419.650000 ;
      RECT 307.500000 418.350000 308.500000 419.650000 ;
      RECT 216.500000 418.350000 299.500000 419.650000 ;
      RECT 207.500000 418.350000 208.500000 419.650000 ;
      RECT 116.500000 418.350000 199.500000 419.650000 ;
      RECT 107.500000 418.350000 108.500000 419.650000 ;
      RECT 66.500000 418.350000 99.500000 419.650000 ;
      RECT 57.500000 418.350000 58.500000 419.650000 ;
      RECT 29.500000 418.350000 49.500000 419.650000 ;
      RECT 15.500000 418.350000 16.500000 419.650000 ;
      RECT 1157.500000 417.650000 1170.500000 418.350000 ;
      RECT 1107.500000 417.650000 1149.500000 418.350000 ;
      RECT 1057.500000 417.650000 1099.500000 418.350000 ;
      RECT 1007.500000 417.650000 1049.500000 418.350000 ;
      RECT 957.500000 417.650000 999.500000 418.350000 ;
      RECT 907.500000 417.650000 949.500000 418.350000 ;
      RECT 857.500000 417.650000 899.500000 418.350000 ;
      RECT 807.500000 417.650000 849.500000 418.350000 ;
      RECT 757.500000 417.650000 799.500000 418.350000 ;
      RECT 707.500000 417.650000 749.500000 418.350000 ;
      RECT 657.500000 417.650000 699.500000 418.350000 ;
      RECT 607.500000 417.650000 649.500000 418.350000 ;
      RECT 557.500000 417.650000 599.500000 418.350000 ;
      RECT 507.500000 417.650000 549.500000 418.350000 ;
      RECT 407.500000 417.650000 499.500000 418.350000 ;
      RECT 357.500000 417.650000 399.500000 418.350000 ;
      RECT 307.500000 417.650000 349.500000 418.350000 ;
      RECT 207.500000 417.650000 299.500000 418.350000 ;
      RECT 107.500000 417.650000 199.500000 418.350000 ;
      RECT 57.500000 417.650000 99.500000 418.350000 ;
      RECT 15.500000 417.650000 49.500000 418.350000 ;
      RECT 1183.500000 416.350000 1186.000000 419.650000 ;
      RECT 1169.500000 416.350000 1170.500000 417.650000 ;
      RECT 1116.500000 416.350000 1149.500000 417.650000 ;
      RECT 1107.500000 416.350000 1108.500000 417.650000 ;
      RECT 1066.500000 416.350000 1099.500000 417.650000 ;
      RECT 1057.500000 416.350000 1058.500000 417.650000 ;
      RECT 1016.500000 416.350000 1049.500000 417.650000 ;
      RECT 1007.500000 416.350000 1008.500000 417.650000 ;
      RECT 966.500000 416.350000 999.500000 417.650000 ;
      RECT 957.500000 416.350000 958.500000 417.650000 ;
      RECT 916.500000 416.350000 949.500000 417.650000 ;
      RECT 907.500000 416.350000 908.500000 417.650000 ;
      RECT 866.500000 416.350000 899.500000 417.650000 ;
      RECT 857.500000 416.350000 858.500000 417.650000 ;
      RECT 816.500000 416.350000 849.500000 417.650000 ;
      RECT 807.500000 416.350000 808.500000 417.650000 ;
      RECT 766.500000 416.350000 799.500000 417.650000 ;
      RECT 757.500000 416.350000 758.500000 417.650000 ;
      RECT 716.500000 416.350000 749.500000 417.650000 ;
      RECT 707.500000 416.350000 708.500000 417.650000 ;
      RECT 666.500000 416.350000 699.500000 417.650000 ;
      RECT 657.500000 416.350000 658.500000 417.650000 ;
      RECT 616.500000 416.350000 649.500000 417.650000 ;
      RECT 607.500000 416.350000 608.500000 417.650000 ;
      RECT 566.500000 416.350000 599.500000 417.650000 ;
      RECT 557.500000 416.350000 558.500000 417.650000 ;
      RECT 516.500000 416.350000 549.500000 417.650000 ;
      RECT 507.500000 416.350000 508.500000 417.650000 ;
      RECT 416.500000 416.350000 499.500000 417.650000 ;
      RECT 407.500000 416.350000 408.500000 417.650000 ;
      RECT 366.500000 416.350000 399.500000 417.650000 ;
      RECT 357.500000 416.350000 358.500000 417.650000 ;
      RECT 316.500000 416.350000 349.500000 417.650000 ;
      RECT 307.500000 416.350000 308.500000 417.650000 ;
      RECT 216.500000 416.350000 299.500000 417.650000 ;
      RECT 207.500000 416.350000 208.500000 417.650000 ;
      RECT 116.500000 416.350000 199.500000 417.650000 ;
      RECT 107.500000 416.350000 108.500000 417.650000 ;
      RECT 66.500000 416.350000 99.500000 417.650000 ;
      RECT 57.500000 416.350000 58.500000 417.650000 ;
      RECT 29.500000 416.350000 49.500000 417.650000 ;
      RECT 15.500000 416.350000 16.500000 417.650000 ;
      RECT 0.000000 416.350000 2.500000 419.650000 ;
      RECT 1169.500000 415.650000 1186.000000 416.350000 ;
      RECT 1116.500000 415.650000 1156.500000 416.350000 ;
      RECT 1066.500000 415.650000 1108.500000 416.350000 ;
      RECT 1016.500000 415.650000 1058.500000 416.350000 ;
      RECT 966.500000 415.650000 1008.500000 416.350000 ;
      RECT 916.500000 415.650000 958.500000 416.350000 ;
      RECT 866.500000 415.650000 908.500000 416.350000 ;
      RECT 816.500000 415.650000 858.500000 416.350000 ;
      RECT 766.500000 415.650000 808.500000 416.350000 ;
      RECT 716.500000 415.650000 758.500000 416.350000 ;
      RECT 666.500000 415.650000 708.500000 416.350000 ;
      RECT 616.500000 415.650000 658.500000 416.350000 ;
      RECT 566.500000 415.650000 608.500000 416.350000 ;
      RECT 516.500000 415.650000 558.500000 416.350000 ;
      RECT 416.500000 415.650000 508.500000 416.350000 ;
      RECT 366.500000 415.650000 408.500000 416.350000 ;
      RECT 316.500000 415.650000 358.500000 416.350000 ;
      RECT 216.500000 415.650000 308.500000 416.350000 ;
      RECT 116.500000 415.650000 208.500000 416.350000 ;
      RECT 66.500000 415.650000 108.500000 416.350000 ;
      RECT 29.500000 415.650000 58.500000 416.350000 ;
      RECT 0.000000 415.650000 16.500000 416.350000 ;
      RECT 1169.500000 414.350000 1170.500000 415.650000 ;
      RECT 1116.500000 414.350000 1149.500000 415.650000 ;
      RECT 1107.500000 414.350000 1108.500000 415.650000 ;
      RECT 1066.500000 414.350000 1099.500000 415.650000 ;
      RECT 1057.500000 414.350000 1058.500000 415.650000 ;
      RECT 1016.500000 414.350000 1049.500000 415.650000 ;
      RECT 1007.500000 414.350000 1008.500000 415.650000 ;
      RECT 966.500000 414.350000 999.500000 415.650000 ;
      RECT 957.500000 414.350000 958.500000 415.650000 ;
      RECT 916.500000 414.350000 949.500000 415.650000 ;
      RECT 907.500000 414.350000 908.500000 415.650000 ;
      RECT 866.500000 414.350000 899.500000 415.650000 ;
      RECT 857.500000 414.350000 858.500000 415.650000 ;
      RECT 816.500000 414.350000 849.500000 415.650000 ;
      RECT 807.500000 414.350000 808.500000 415.650000 ;
      RECT 766.500000 414.350000 799.500000 415.650000 ;
      RECT 757.500000 414.350000 758.500000 415.650000 ;
      RECT 716.500000 414.350000 749.500000 415.650000 ;
      RECT 707.500000 414.350000 708.500000 415.650000 ;
      RECT 666.500000 414.350000 699.500000 415.650000 ;
      RECT 657.500000 414.350000 658.500000 415.650000 ;
      RECT 616.500000 414.350000 649.500000 415.650000 ;
      RECT 607.500000 414.350000 608.500000 415.650000 ;
      RECT 566.500000 414.350000 599.500000 415.650000 ;
      RECT 557.500000 414.350000 558.500000 415.650000 ;
      RECT 516.500000 414.350000 549.500000 415.650000 ;
      RECT 507.500000 414.350000 508.500000 415.650000 ;
      RECT 416.500000 414.350000 499.500000 415.650000 ;
      RECT 407.500000 414.350000 408.500000 415.650000 ;
      RECT 366.500000 414.350000 399.500000 415.650000 ;
      RECT 357.500000 414.350000 358.500000 415.650000 ;
      RECT 316.500000 414.350000 349.500000 415.650000 ;
      RECT 307.500000 414.350000 308.500000 415.650000 ;
      RECT 216.500000 414.350000 299.500000 415.650000 ;
      RECT 207.500000 414.350000 208.500000 415.650000 ;
      RECT 116.500000 414.350000 199.500000 415.650000 ;
      RECT 107.500000 414.350000 108.500000 415.650000 ;
      RECT 66.500000 414.350000 99.500000 415.650000 ;
      RECT 57.500000 414.350000 58.500000 415.650000 ;
      RECT 29.500000 414.350000 49.500000 415.650000 ;
      RECT 15.500000 414.350000 16.500000 415.650000 ;
      RECT 1157.500000 413.650000 1170.500000 414.350000 ;
      RECT 1107.500000 413.650000 1149.500000 414.350000 ;
      RECT 1057.500000 413.650000 1099.500000 414.350000 ;
      RECT 1007.500000 413.650000 1049.500000 414.350000 ;
      RECT 957.500000 413.650000 999.500000 414.350000 ;
      RECT 907.500000 413.650000 949.500000 414.350000 ;
      RECT 857.500000 413.650000 899.500000 414.350000 ;
      RECT 807.500000 413.650000 849.500000 414.350000 ;
      RECT 757.500000 413.650000 799.500000 414.350000 ;
      RECT 707.500000 413.650000 749.500000 414.350000 ;
      RECT 657.500000 413.650000 699.500000 414.350000 ;
      RECT 607.500000 413.650000 649.500000 414.350000 ;
      RECT 557.500000 413.650000 599.500000 414.350000 ;
      RECT 507.500000 413.650000 549.500000 414.350000 ;
      RECT 407.500000 413.650000 499.500000 414.350000 ;
      RECT 357.500000 413.650000 399.500000 414.350000 ;
      RECT 307.500000 413.650000 349.500000 414.350000 ;
      RECT 207.500000 413.650000 299.500000 414.350000 ;
      RECT 107.500000 413.650000 199.500000 414.350000 ;
      RECT 57.500000 413.650000 99.500000 414.350000 ;
      RECT 15.500000 413.650000 49.500000 414.350000 ;
      RECT 1183.500000 412.350000 1186.000000 415.650000 ;
      RECT 1169.500000 412.350000 1170.500000 413.650000 ;
      RECT 1116.500000 412.350000 1149.500000 413.650000 ;
      RECT 1107.500000 412.350000 1108.500000 413.650000 ;
      RECT 1066.500000 412.350000 1099.500000 413.650000 ;
      RECT 1057.500000 412.350000 1058.500000 413.650000 ;
      RECT 1016.500000 412.350000 1049.500000 413.650000 ;
      RECT 1007.500000 412.350000 1008.500000 413.650000 ;
      RECT 966.500000 412.350000 999.500000 413.650000 ;
      RECT 957.500000 412.350000 958.500000 413.650000 ;
      RECT 916.500000 412.350000 949.500000 413.650000 ;
      RECT 907.500000 412.350000 908.500000 413.650000 ;
      RECT 866.500000 412.350000 899.500000 413.650000 ;
      RECT 857.500000 412.350000 858.500000 413.650000 ;
      RECT 816.500000 412.350000 849.500000 413.650000 ;
      RECT 807.500000 412.350000 808.500000 413.650000 ;
      RECT 766.500000 412.350000 799.500000 413.650000 ;
      RECT 757.500000 412.350000 758.500000 413.650000 ;
      RECT 716.500000 412.350000 749.500000 413.650000 ;
      RECT 707.500000 412.350000 708.500000 413.650000 ;
      RECT 666.500000 412.350000 699.500000 413.650000 ;
      RECT 657.500000 412.350000 658.500000 413.650000 ;
      RECT 616.500000 412.350000 649.500000 413.650000 ;
      RECT 607.500000 412.350000 608.500000 413.650000 ;
      RECT 566.500000 412.350000 599.500000 413.650000 ;
      RECT 557.500000 412.350000 558.500000 413.650000 ;
      RECT 516.500000 412.350000 549.500000 413.650000 ;
      RECT 507.500000 412.350000 508.500000 413.650000 ;
      RECT 416.500000 412.350000 499.500000 413.650000 ;
      RECT 407.500000 412.350000 408.500000 413.650000 ;
      RECT 366.500000 412.350000 399.500000 413.650000 ;
      RECT 357.500000 412.350000 358.500000 413.650000 ;
      RECT 316.500000 412.350000 349.500000 413.650000 ;
      RECT 307.500000 412.350000 308.500000 413.650000 ;
      RECT 216.500000 412.350000 299.500000 413.650000 ;
      RECT 207.500000 412.350000 208.500000 413.650000 ;
      RECT 116.500000 412.350000 199.500000 413.650000 ;
      RECT 107.500000 412.350000 108.500000 413.650000 ;
      RECT 66.500000 412.350000 99.500000 413.650000 ;
      RECT 57.500000 412.350000 58.500000 413.650000 ;
      RECT 29.500000 412.350000 49.500000 413.650000 ;
      RECT 15.500000 412.350000 16.500000 413.650000 ;
      RECT 0.000000 412.350000 2.500000 415.650000 ;
      RECT 1169.500000 411.650000 1186.000000 412.350000 ;
      RECT 1116.500000 411.650000 1156.500000 412.350000 ;
      RECT 1066.500000 411.650000 1108.500000 412.350000 ;
      RECT 1016.500000 411.650000 1058.500000 412.350000 ;
      RECT 966.500000 411.650000 1008.500000 412.350000 ;
      RECT 916.500000 411.650000 958.500000 412.350000 ;
      RECT 866.500000 411.650000 908.500000 412.350000 ;
      RECT 816.500000 411.650000 858.500000 412.350000 ;
      RECT 766.500000 411.650000 808.500000 412.350000 ;
      RECT 716.500000 411.650000 758.500000 412.350000 ;
      RECT 666.500000 411.650000 708.500000 412.350000 ;
      RECT 616.500000 411.650000 658.500000 412.350000 ;
      RECT 566.500000 411.650000 608.500000 412.350000 ;
      RECT 516.500000 411.650000 558.500000 412.350000 ;
      RECT 416.500000 411.650000 508.500000 412.350000 ;
      RECT 366.500000 411.650000 408.500000 412.350000 ;
      RECT 316.500000 411.650000 358.500000 412.350000 ;
      RECT 216.500000 411.650000 308.500000 412.350000 ;
      RECT 116.500000 411.650000 208.500000 412.350000 ;
      RECT 66.500000 411.650000 108.500000 412.350000 ;
      RECT 29.500000 411.650000 58.500000 412.350000 ;
      RECT 0.000000 411.650000 16.500000 412.350000 ;
      RECT 1169.500000 410.350000 1170.500000 411.650000 ;
      RECT 1116.500000 410.350000 1149.500000 411.650000 ;
      RECT 1107.500000 410.350000 1108.500000 411.650000 ;
      RECT 1066.500000 410.350000 1099.500000 411.650000 ;
      RECT 1057.500000 410.350000 1058.500000 411.650000 ;
      RECT 1016.500000 410.350000 1049.500000 411.650000 ;
      RECT 1007.500000 410.350000 1008.500000 411.650000 ;
      RECT 966.500000 410.350000 999.500000 411.650000 ;
      RECT 957.500000 410.350000 958.500000 411.650000 ;
      RECT 916.500000 410.350000 949.500000 411.650000 ;
      RECT 907.500000 410.350000 908.500000 411.650000 ;
      RECT 866.500000 410.350000 899.500000 411.650000 ;
      RECT 857.500000 410.350000 858.500000 411.650000 ;
      RECT 816.500000 410.350000 849.500000 411.650000 ;
      RECT 807.500000 410.350000 808.500000 411.650000 ;
      RECT 766.500000 410.350000 799.500000 411.650000 ;
      RECT 757.500000 410.350000 758.500000 411.650000 ;
      RECT 716.500000 410.350000 749.500000 411.650000 ;
      RECT 707.500000 410.350000 708.500000 411.650000 ;
      RECT 666.500000 410.350000 699.500000 411.650000 ;
      RECT 657.500000 410.350000 658.500000 411.650000 ;
      RECT 616.500000 410.350000 649.500000 411.650000 ;
      RECT 607.500000 410.350000 608.500000 411.650000 ;
      RECT 566.500000 410.350000 599.500000 411.650000 ;
      RECT 557.500000 410.350000 558.500000 411.650000 ;
      RECT 516.500000 410.350000 549.500000 411.650000 ;
      RECT 507.500000 410.350000 508.500000 411.650000 ;
      RECT 416.500000 410.350000 499.500000 411.650000 ;
      RECT 407.500000 410.350000 408.500000 411.650000 ;
      RECT 366.500000 410.350000 399.500000 411.650000 ;
      RECT 357.500000 410.350000 358.500000 411.650000 ;
      RECT 316.500000 410.350000 349.500000 411.650000 ;
      RECT 307.500000 410.350000 308.500000 411.650000 ;
      RECT 216.500000 410.350000 299.500000 411.650000 ;
      RECT 207.500000 410.350000 208.500000 411.650000 ;
      RECT 116.500000 410.350000 199.500000 411.650000 ;
      RECT 107.500000 410.350000 108.500000 411.650000 ;
      RECT 66.500000 410.350000 99.500000 411.650000 ;
      RECT 57.500000 410.350000 58.500000 411.650000 ;
      RECT 29.500000 410.350000 49.500000 411.650000 ;
      RECT 15.500000 410.350000 16.500000 411.650000 ;
      RECT 1157.500000 409.650000 1170.500000 410.350000 ;
      RECT 1107.500000 409.650000 1149.500000 410.350000 ;
      RECT 1057.500000 409.650000 1099.500000 410.350000 ;
      RECT 1007.500000 409.650000 1049.500000 410.350000 ;
      RECT 957.500000 409.650000 999.500000 410.350000 ;
      RECT 907.500000 409.650000 949.500000 410.350000 ;
      RECT 857.500000 409.650000 899.500000 410.350000 ;
      RECT 807.500000 409.650000 849.500000 410.350000 ;
      RECT 757.500000 409.650000 799.500000 410.350000 ;
      RECT 707.500000 409.650000 749.500000 410.350000 ;
      RECT 657.500000 409.650000 699.500000 410.350000 ;
      RECT 607.500000 409.650000 649.500000 410.350000 ;
      RECT 557.500000 409.650000 599.500000 410.350000 ;
      RECT 507.500000 409.650000 549.500000 410.350000 ;
      RECT 407.500000 409.650000 499.500000 410.350000 ;
      RECT 357.500000 409.650000 399.500000 410.350000 ;
      RECT 307.500000 409.650000 349.500000 410.350000 ;
      RECT 207.500000 409.650000 299.500000 410.350000 ;
      RECT 107.500000 409.650000 199.500000 410.350000 ;
      RECT 57.500000 409.650000 99.500000 410.350000 ;
      RECT 15.500000 409.650000 49.500000 410.350000 ;
      RECT 1183.500000 408.350000 1186.000000 411.650000 ;
      RECT 1169.500000 408.350000 1170.500000 409.650000 ;
      RECT 1116.500000 408.350000 1149.500000 409.650000 ;
      RECT 1107.500000 408.350000 1108.500000 409.650000 ;
      RECT 1066.500000 408.350000 1099.500000 409.650000 ;
      RECT 1057.500000 408.350000 1058.500000 409.650000 ;
      RECT 1016.500000 408.350000 1049.500000 409.650000 ;
      RECT 1007.500000 408.350000 1008.500000 409.650000 ;
      RECT 966.500000 408.350000 999.500000 409.650000 ;
      RECT 957.500000 408.350000 958.500000 409.650000 ;
      RECT 916.500000 408.350000 949.500000 409.650000 ;
      RECT 907.500000 408.350000 908.500000 409.650000 ;
      RECT 866.500000 408.350000 899.500000 409.650000 ;
      RECT 857.500000 408.350000 858.500000 409.650000 ;
      RECT 816.500000 408.350000 849.500000 409.650000 ;
      RECT 807.500000 408.350000 808.500000 409.650000 ;
      RECT 766.500000 408.350000 799.500000 409.650000 ;
      RECT 757.500000 408.350000 758.500000 409.650000 ;
      RECT 716.500000 408.350000 749.500000 409.650000 ;
      RECT 707.500000 408.350000 708.500000 409.650000 ;
      RECT 666.500000 408.350000 699.500000 409.650000 ;
      RECT 657.500000 408.350000 658.500000 409.650000 ;
      RECT 616.500000 408.350000 649.500000 409.650000 ;
      RECT 607.500000 408.350000 608.500000 409.650000 ;
      RECT 566.500000 408.350000 599.500000 409.650000 ;
      RECT 557.500000 408.350000 558.500000 409.650000 ;
      RECT 516.500000 408.350000 549.500000 409.650000 ;
      RECT 507.500000 408.350000 508.500000 409.650000 ;
      RECT 416.500000 408.350000 499.500000 409.650000 ;
      RECT 407.500000 408.350000 408.500000 409.650000 ;
      RECT 366.500000 408.350000 399.500000 409.650000 ;
      RECT 357.500000 408.350000 358.500000 409.650000 ;
      RECT 316.500000 408.350000 349.500000 409.650000 ;
      RECT 307.500000 408.350000 308.500000 409.650000 ;
      RECT 216.500000 408.350000 299.500000 409.650000 ;
      RECT 207.500000 408.350000 208.500000 409.650000 ;
      RECT 116.500000 408.350000 199.500000 409.650000 ;
      RECT 107.500000 408.350000 108.500000 409.650000 ;
      RECT 66.500000 408.350000 99.500000 409.650000 ;
      RECT 57.500000 408.350000 58.500000 409.650000 ;
      RECT 29.500000 408.350000 49.500000 409.650000 ;
      RECT 15.500000 408.350000 16.500000 409.650000 ;
      RECT 0.000000 408.350000 2.500000 411.650000 ;
      RECT 1169.500000 407.650000 1186.000000 408.350000 ;
      RECT 1116.500000 407.650000 1156.500000 408.350000 ;
      RECT 1066.500000 407.650000 1108.500000 408.350000 ;
      RECT 1016.500000 407.650000 1058.500000 408.350000 ;
      RECT 966.500000 407.650000 1008.500000 408.350000 ;
      RECT 916.500000 407.650000 958.500000 408.350000 ;
      RECT 866.500000 407.650000 908.500000 408.350000 ;
      RECT 816.500000 407.650000 858.500000 408.350000 ;
      RECT 766.500000 407.650000 808.500000 408.350000 ;
      RECT 716.500000 407.650000 758.500000 408.350000 ;
      RECT 666.500000 407.650000 708.500000 408.350000 ;
      RECT 616.500000 407.650000 658.500000 408.350000 ;
      RECT 566.500000 407.650000 608.500000 408.350000 ;
      RECT 516.500000 407.650000 558.500000 408.350000 ;
      RECT 416.500000 407.650000 508.500000 408.350000 ;
      RECT 366.500000 407.650000 408.500000 408.350000 ;
      RECT 316.500000 407.650000 358.500000 408.350000 ;
      RECT 216.500000 407.650000 308.500000 408.350000 ;
      RECT 116.500000 407.650000 208.500000 408.350000 ;
      RECT 66.500000 407.650000 108.500000 408.350000 ;
      RECT 29.500000 407.650000 58.500000 408.350000 ;
      RECT 0.000000 407.650000 16.500000 408.350000 ;
      RECT 1169.500000 406.350000 1170.500000 407.650000 ;
      RECT 1116.500000 406.350000 1149.500000 407.650000 ;
      RECT 1107.500000 406.350000 1108.500000 407.650000 ;
      RECT 1066.500000 406.350000 1099.500000 407.650000 ;
      RECT 1057.500000 406.350000 1058.500000 407.650000 ;
      RECT 1016.500000 406.350000 1049.500000 407.650000 ;
      RECT 1007.500000 406.350000 1008.500000 407.650000 ;
      RECT 966.500000 406.350000 999.500000 407.650000 ;
      RECT 957.500000 406.350000 958.500000 407.650000 ;
      RECT 916.500000 406.350000 949.500000 407.650000 ;
      RECT 907.500000 406.350000 908.500000 407.650000 ;
      RECT 866.500000 406.350000 899.500000 407.650000 ;
      RECT 857.500000 406.350000 858.500000 407.650000 ;
      RECT 816.500000 406.350000 849.500000 407.650000 ;
      RECT 807.500000 406.350000 808.500000 407.650000 ;
      RECT 766.500000 406.350000 799.500000 407.650000 ;
      RECT 757.500000 406.350000 758.500000 407.650000 ;
      RECT 716.500000 406.350000 749.500000 407.650000 ;
      RECT 707.500000 406.350000 708.500000 407.650000 ;
      RECT 666.500000 406.350000 699.500000 407.650000 ;
      RECT 657.500000 406.350000 658.500000 407.650000 ;
      RECT 616.500000 406.350000 649.500000 407.650000 ;
      RECT 607.500000 406.350000 608.500000 407.650000 ;
      RECT 566.500000 406.350000 599.500000 407.650000 ;
      RECT 557.500000 406.350000 558.500000 407.650000 ;
      RECT 516.500000 406.350000 549.500000 407.650000 ;
      RECT 507.500000 406.350000 508.500000 407.650000 ;
      RECT 416.500000 406.350000 499.500000 407.650000 ;
      RECT 407.500000 406.350000 408.500000 407.650000 ;
      RECT 366.500000 406.350000 399.500000 407.650000 ;
      RECT 357.500000 406.350000 358.500000 407.650000 ;
      RECT 316.500000 406.350000 349.500000 407.650000 ;
      RECT 307.500000 406.350000 308.500000 407.650000 ;
      RECT 216.500000 406.350000 299.500000 407.650000 ;
      RECT 207.500000 406.350000 208.500000 407.650000 ;
      RECT 116.500000 406.350000 199.500000 407.650000 ;
      RECT 107.500000 406.350000 108.500000 407.650000 ;
      RECT 66.500000 406.350000 99.500000 407.650000 ;
      RECT 57.500000 406.350000 58.500000 407.650000 ;
      RECT 29.500000 406.350000 49.500000 407.650000 ;
      RECT 15.500000 406.350000 16.500000 407.650000 ;
      RECT 1157.500000 405.650000 1170.500000 406.350000 ;
      RECT 1107.500000 405.650000 1149.500000 406.350000 ;
      RECT 1057.500000 405.650000 1099.500000 406.350000 ;
      RECT 1007.500000 405.650000 1049.500000 406.350000 ;
      RECT 957.500000 405.650000 999.500000 406.350000 ;
      RECT 907.500000 405.650000 949.500000 406.350000 ;
      RECT 857.500000 405.650000 899.500000 406.350000 ;
      RECT 807.500000 405.650000 849.500000 406.350000 ;
      RECT 757.500000 405.650000 799.500000 406.350000 ;
      RECT 707.500000 405.650000 749.500000 406.350000 ;
      RECT 657.500000 405.650000 699.500000 406.350000 ;
      RECT 607.500000 405.650000 649.500000 406.350000 ;
      RECT 557.500000 405.650000 599.500000 406.350000 ;
      RECT 507.500000 405.650000 549.500000 406.350000 ;
      RECT 407.500000 405.650000 499.500000 406.350000 ;
      RECT 357.500000 405.650000 399.500000 406.350000 ;
      RECT 307.500000 405.650000 349.500000 406.350000 ;
      RECT 207.500000 405.650000 299.500000 406.350000 ;
      RECT 107.500000 405.650000 199.500000 406.350000 ;
      RECT 57.500000 405.650000 99.500000 406.350000 ;
      RECT 15.500000 405.650000 49.500000 406.350000 ;
      RECT 1183.500000 404.350000 1186.000000 407.650000 ;
      RECT 1169.500000 404.350000 1170.500000 405.650000 ;
      RECT 1116.500000 404.350000 1149.500000 405.650000 ;
      RECT 1107.500000 404.350000 1108.500000 405.650000 ;
      RECT 1066.500000 404.350000 1099.500000 405.650000 ;
      RECT 1057.500000 404.350000 1058.500000 405.650000 ;
      RECT 1016.500000 404.350000 1049.500000 405.650000 ;
      RECT 1007.500000 404.350000 1008.500000 405.650000 ;
      RECT 966.500000 404.350000 999.500000 405.650000 ;
      RECT 957.500000 404.350000 958.500000 405.650000 ;
      RECT 916.500000 404.350000 949.500000 405.650000 ;
      RECT 907.500000 404.350000 908.500000 405.650000 ;
      RECT 866.500000 404.350000 899.500000 405.650000 ;
      RECT 857.500000 404.350000 858.500000 405.650000 ;
      RECT 816.500000 404.350000 849.500000 405.650000 ;
      RECT 807.500000 404.350000 808.500000 405.650000 ;
      RECT 766.500000 404.350000 799.500000 405.650000 ;
      RECT 757.500000 404.350000 758.500000 405.650000 ;
      RECT 716.500000 404.350000 749.500000 405.650000 ;
      RECT 707.500000 404.350000 708.500000 405.650000 ;
      RECT 666.500000 404.350000 699.500000 405.650000 ;
      RECT 657.500000 404.350000 658.500000 405.650000 ;
      RECT 616.500000 404.350000 649.500000 405.650000 ;
      RECT 607.500000 404.350000 608.500000 405.650000 ;
      RECT 566.500000 404.350000 599.500000 405.650000 ;
      RECT 557.500000 404.350000 558.500000 405.650000 ;
      RECT 516.500000 404.350000 549.500000 405.650000 ;
      RECT 507.500000 404.350000 508.500000 405.650000 ;
      RECT 416.500000 404.350000 499.500000 405.650000 ;
      RECT 407.500000 404.350000 408.500000 405.650000 ;
      RECT 366.500000 404.350000 399.500000 405.650000 ;
      RECT 357.500000 404.350000 358.500000 405.650000 ;
      RECT 316.500000 404.350000 349.500000 405.650000 ;
      RECT 307.500000 404.350000 308.500000 405.650000 ;
      RECT 216.500000 404.350000 299.500000 405.650000 ;
      RECT 207.500000 404.350000 208.500000 405.650000 ;
      RECT 116.500000 404.350000 199.500000 405.650000 ;
      RECT 107.500000 404.350000 108.500000 405.650000 ;
      RECT 66.500000 404.350000 99.500000 405.650000 ;
      RECT 57.500000 404.350000 58.500000 405.650000 ;
      RECT 29.500000 404.350000 49.500000 405.650000 ;
      RECT 15.500000 404.350000 16.500000 405.650000 ;
      RECT 0.000000 404.350000 2.500000 407.650000 ;
      RECT 1169.500000 403.650000 1186.000000 404.350000 ;
      RECT 1116.500000 403.650000 1156.500000 404.350000 ;
      RECT 1066.500000 403.650000 1108.500000 404.350000 ;
      RECT 1016.500000 403.650000 1058.500000 404.350000 ;
      RECT 966.500000 403.650000 1008.500000 404.350000 ;
      RECT 916.500000 403.650000 958.500000 404.350000 ;
      RECT 866.500000 403.650000 908.500000 404.350000 ;
      RECT 816.500000 403.650000 858.500000 404.350000 ;
      RECT 766.500000 403.650000 808.500000 404.350000 ;
      RECT 716.500000 403.650000 758.500000 404.350000 ;
      RECT 666.500000 403.650000 708.500000 404.350000 ;
      RECT 616.500000 403.650000 658.500000 404.350000 ;
      RECT 566.500000 403.650000 608.500000 404.350000 ;
      RECT 516.500000 403.650000 558.500000 404.350000 ;
      RECT 416.500000 403.650000 508.500000 404.350000 ;
      RECT 366.500000 403.650000 408.500000 404.350000 ;
      RECT 316.500000 403.650000 358.500000 404.350000 ;
      RECT 216.500000 403.650000 308.500000 404.350000 ;
      RECT 116.500000 403.650000 208.500000 404.350000 ;
      RECT 66.500000 403.650000 108.500000 404.350000 ;
      RECT 29.500000 403.650000 58.500000 404.350000 ;
      RECT 0.000000 403.650000 16.500000 404.350000 ;
      RECT 1169.500000 402.350000 1170.500000 403.650000 ;
      RECT 1116.500000 402.350000 1149.500000 403.650000 ;
      RECT 1107.500000 402.350000 1108.500000 403.650000 ;
      RECT 1066.500000 402.350000 1099.500000 403.650000 ;
      RECT 1057.500000 402.350000 1058.500000 403.650000 ;
      RECT 1016.500000 402.350000 1049.500000 403.650000 ;
      RECT 1007.500000 402.350000 1008.500000 403.650000 ;
      RECT 966.500000 402.350000 999.500000 403.650000 ;
      RECT 957.500000 402.350000 958.500000 403.650000 ;
      RECT 916.500000 402.350000 949.500000 403.650000 ;
      RECT 907.500000 402.350000 908.500000 403.650000 ;
      RECT 866.500000 402.350000 899.500000 403.650000 ;
      RECT 857.500000 402.350000 858.500000 403.650000 ;
      RECT 816.500000 402.350000 849.500000 403.650000 ;
      RECT 807.500000 402.350000 808.500000 403.650000 ;
      RECT 766.500000 402.350000 799.500000 403.650000 ;
      RECT 757.500000 402.350000 758.500000 403.650000 ;
      RECT 716.500000 402.350000 749.500000 403.650000 ;
      RECT 707.500000 402.350000 708.500000 403.650000 ;
      RECT 666.500000 402.350000 699.500000 403.650000 ;
      RECT 657.500000 402.350000 658.500000 403.650000 ;
      RECT 616.500000 402.350000 649.500000 403.650000 ;
      RECT 607.500000 402.350000 608.500000 403.650000 ;
      RECT 566.500000 402.350000 599.500000 403.650000 ;
      RECT 557.500000 402.350000 558.500000 403.650000 ;
      RECT 516.500000 402.350000 549.500000 403.650000 ;
      RECT 507.500000 402.350000 508.500000 403.650000 ;
      RECT 416.500000 402.350000 499.500000 403.650000 ;
      RECT 407.500000 402.350000 408.500000 403.650000 ;
      RECT 366.500000 402.350000 399.500000 403.650000 ;
      RECT 357.500000 402.350000 358.500000 403.650000 ;
      RECT 316.500000 402.350000 349.500000 403.650000 ;
      RECT 307.500000 402.350000 308.500000 403.650000 ;
      RECT 216.500000 402.350000 249.500000 403.650000 ;
      RECT 207.500000 402.350000 208.500000 403.650000 ;
      RECT 116.500000 402.350000 149.500000 403.650000 ;
      RECT 107.500000 402.350000 108.500000 403.650000 ;
      RECT 66.500000 402.350000 99.500000 403.650000 ;
      RECT 57.500000 402.350000 58.500000 403.650000 ;
      RECT 29.500000 402.350000 49.500000 403.650000 ;
      RECT 15.500000 402.350000 16.500000 403.650000 ;
      RECT 1157.500000 401.650000 1170.500000 402.350000 ;
      RECT 1107.500000 401.650000 1149.500000 402.350000 ;
      RECT 1057.500000 401.650000 1099.500000 402.350000 ;
      RECT 1007.500000 401.650000 1049.500000 402.350000 ;
      RECT 957.500000 401.650000 999.500000 402.350000 ;
      RECT 907.500000 401.650000 949.500000 402.350000 ;
      RECT 857.500000 401.650000 899.500000 402.350000 ;
      RECT 807.500000 401.650000 849.500000 402.350000 ;
      RECT 757.500000 401.650000 799.500000 402.350000 ;
      RECT 707.500000 401.650000 749.500000 402.350000 ;
      RECT 657.500000 401.650000 699.500000 402.350000 ;
      RECT 607.500000 401.650000 649.500000 402.350000 ;
      RECT 557.500000 401.650000 599.500000 402.350000 ;
      RECT 507.500000 401.650000 549.500000 402.350000 ;
      RECT 407.500000 401.650000 499.500000 402.350000 ;
      RECT 357.500000 401.650000 399.500000 402.350000 ;
      RECT 307.500000 401.650000 349.500000 402.350000 ;
      RECT 257.500000 401.650000 299.500000 403.650000 ;
      RECT 207.500000 401.650000 249.500000 402.350000 ;
      RECT 157.500000 401.650000 199.500000 403.650000 ;
      RECT 107.500000 401.650000 149.500000 402.350000 ;
      RECT 57.500000 401.650000 99.500000 402.350000 ;
      RECT 15.500000 401.650000 49.500000 402.350000 ;
      RECT 1183.500000 400.350000 1186.000000 403.650000 ;
      RECT 1169.500000 400.350000 1170.500000 401.650000 ;
      RECT 1116.500000 400.350000 1149.500000 401.650000 ;
      RECT 1107.500000 400.350000 1108.500000 401.650000 ;
      RECT 1066.500000 400.350000 1099.500000 401.650000 ;
      RECT 1057.500000 400.350000 1058.500000 401.650000 ;
      RECT 1016.500000 400.350000 1049.500000 401.650000 ;
      RECT 1007.500000 400.350000 1008.500000 401.650000 ;
      RECT 966.500000 400.350000 999.500000 401.650000 ;
      RECT 957.500000 400.350000 958.500000 401.650000 ;
      RECT 916.500000 400.350000 949.500000 401.650000 ;
      RECT 907.500000 400.350000 908.500000 401.650000 ;
      RECT 866.500000 400.350000 899.500000 401.650000 ;
      RECT 857.500000 400.350000 858.500000 401.650000 ;
      RECT 816.500000 400.350000 849.500000 401.650000 ;
      RECT 807.500000 400.350000 808.500000 401.650000 ;
      RECT 766.500000 400.350000 799.500000 401.650000 ;
      RECT 757.500000 400.350000 758.500000 401.650000 ;
      RECT 716.500000 400.350000 749.500000 401.650000 ;
      RECT 707.500000 400.350000 708.500000 401.650000 ;
      RECT 666.500000 400.350000 699.500000 401.650000 ;
      RECT 657.500000 400.350000 658.500000 401.650000 ;
      RECT 616.500000 400.350000 649.500000 401.650000 ;
      RECT 607.500000 400.350000 608.500000 401.650000 ;
      RECT 566.500000 400.350000 599.500000 401.650000 ;
      RECT 557.500000 400.350000 558.500000 401.650000 ;
      RECT 516.500000 400.350000 549.500000 401.650000 ;
      RECT 507.500000 400.350000 508.500000 401.650000 ;
      RECT 416.500000 400.350000 499.500000 401.650000 ;
      RECT 407.500000 400.350000 408.500000 401.650000 ;
      RECT 366.500000 400.350000 399.500000 401.650000 ;
      RECT 357.500000 400.350000 358.500000 401.650000 ;
      RECT 316.500000 400.350000 349.500000 401.650000 ;
      RECT 307.500000 400.350000 308.500000 401.650000 ;
      RECT 266.500000 400.350000 299.500000 401.650000 ;
      RECT 257.500000 400.350000 258.500000 401.650000 ;
      RECT 216.500000 400.350000 249.500000 401.650000 ;
      RECT 207.500000 400.350000 208.500000 401.650000 ;
      RECT 166.500000 400.350000 199.500000 401.650000 ;
      RECT 157.500000 400.350000 158.500000 401.650000 ;
      RECT 116.500000 400.350000 149.500000 401.650000 ;
      RECT 107.500000 400.350000 108.500000 401.650000 ;
      RECT 66.500000 400.350000 99.500000 401.650000 ;
      RECT 57.500000 400.350000 58.500000 401.650000 ;
      RECT 29.500000 400.350000 49.500000 401.650000 ;
      RECT 15.500000 400.350000 16.500000 401.650000 ;
      RECT 0.000000 400.350000 2.500000 403.650000 ;
      RECT 1169.500000 399.650000 1186.000000 400.350000 ;
      RECT 1116.500000 399.650000 1156.500000 400.350000 ;
      RECT 1066.500000 399.650000 1108.500000 400.350000 ;
      RECT 1016.500000 399.650000 1058.500000 400.350000 ;
      RECT 966.500000 399.650000 1008.500000 400.350000 ;
      RECT 916.500000 399.650000 958.500000 400.350000 ;
      RECT 866.500000 399.650000 908.500000 400.350000 ;
      RECT 816.500000 399.650000 858.500000 400.350000 ;
      RECT 766.500000 399.650000 808.500000 400.350000 ;
      RECT 716.500000 399.650000 758.500000 400.350000 ;
      RECT 666.500000 399.650000 708.500000 400.350000 ;
      RECT 616.500000 399.650000 658.500000 400.350000 ;
      RECT 566.500000 399.650000 608.500000 400.350000 ;
      RECT 516.500000 399.650000 558.500000 400.350000 ;
      RECT 416.500000 399.650000 508.500000 400.350000 ;
      RECT 366.500000 399.650000 408.500000 400.350000 ;
      RECT 316.500000 399.650000 358.500000 400.350000 ;
      RECT 266.500000 399.650000 308.500000 400.350000 ;
      RECT 216.500000 399.650000 258.500000 400.350000 ;
      RECT 166.500000 399.650000 208.500000 400.350000 ;
      RECT 116.500000 399.650000 158.500000 400.350000 ;
      RECT 66.500000 399.650000 108.500000 400.350000 ;
      RECT 29.500000 399.650000 58.500000 400.350000 ;
      RECT 0.000000 399.650000 16.500000 400.350000 ;
      RECT 0.000000 399.170000 2.500000 399.650000 ;
      RECT 1183.500000 399.165000 1186.000000 399.650000 ;
      RECT 1169.500000 398.350000 1170.500000 399.650000 ;
      RECT 1116.500000 398.350000 1149.500000 399.650000 ;
      RECT 1107.500000 398.350000 1108.500000 399.650000 ;
      RECT 1066.500000 398.350000 1099.500000 399.650000 ;
      RECT 1057.500000 398.350000 1058.500000 399.650000 ;
      RECT 1016.500000 398.350000 1049.500000 399.650000 ;
      RECT 1007.500000 398.350000 1008.500000 399.650000 ;
      RECT 966.500000 398.350000 999.500000 399.650000 ;
      RECT 957.500000 398.350000 958.500000 399.650000 ;
      RECT 916.500000 398.350000 949.500000 399.650000 ;
      RECT 907.500000 398.350000 908.500000 399.650000 ;
      RECT 866.500000 398.350000 899.500000 399.650000 ;
      RECT 857.500000 398.350000 858.500000 399.650000 ;
      RECT 816.500000 398.350000 849.500000 399.650000 ;
      RECT 807.500000 398.350000 808.500000 399.650000 ;
      RECT 766.500000 398.350000 799.500000 399.650000 ;
      RECT 757.500000 398.350000 758.500000 399.650000 ;
      RECT 716.500000 398.350000 749.500000 399.650000 ;
      RECT 707.500000 398.350000 708.500000 399.650000 ;
      RECT 666.500000 398.350000 699.500000 399.650000 ;
      RECT 657.500000 398.350000 658.500000 399.650000 ;
      RECT 616.500000 398.350000 649.500000 399.650000 ;
      RECT 607.500000 398.350000 608.500000 399.650000 ;
      RECT 566.500000 398.350000 599.500000 399.650000 ;
      RECT 557.500000 398.350000 558.500000 399.650000 ;
      RECT 516.500000 398.350000 549.500000 399.650000 ;
      RECT 507.500000 398.350000 508.500000 399.650000 ;
      RECT 416.500000 398.350000 449.500000 399.650000 ;
      RECT 407.500000 398.350000 408.500000 399.650000 ;
      RECT 366.500000 398.350000 399.500000 399.650000 ;
      RECT 357.500000 398.350000 358.500000 399.650000 ;
      RECT 316.500000 398.350000 349.500000 399.650000 ;
      RECT 307.500000 398.350000 308.500000 399.650000 ;
      RECT 266.500000 398.350000 299.500000 399.650000 ;
      RECT 257.500000 398.350000 258.500000 399.650000 ;
      RECT 216.500000 398.350000 249.500000 399.650000 ;
      RECT 207.500000 398.350000 208.500000 399.650000 ;
      RECT 166.500000 398.350000 199.500000 399.650000 ;
      RECT 157.500000 398.350000 158.500000 399.650000 ;
      RECT 116.500000 398.350000 149.500000 399.650000 ;
      RECT 107.500000 398.350000 108.500000 399.650000 ;
      RECT 66.500000 398.350000 99.500000 399.650000 ;
      RECT 57.500000 398.350000 58.500000 399.650000 ;
      RECT 29.500000 398.350000 49.500000 399.650000 ;
      RECT 15.500000 398.350000 16.500000 399.650000 ;
      RECT 1157.500000 397.650000 1170.500000 398.350000 ;
      RECT 1107.500000 397.650000 1149.500000 398.350000 ;
      RECT 1057.500000 397.650000 1099.500000 398.350000 ;
      RECT 1007.500000 397.650000 1049.500000 398.350000 ;
      RECT 957.500000 397.650000 999.500000 398.350000 ;
      RECT 907.500000 397.650000 949.500000 398.350000 ;
      RECT 857.500000 397.650000 899.500000 398.350000 ;
      RECT 807.500000 397.650000 849.500000 398.350000 ;
      RECT 757.500000 397.650000 799.500000 398.350000 ;
      RECT 707.500000 397.650000 749.500000 398.350000 ;
      RECT 657.500000 397.650000 699.500000 398.350000 ;
      RECT 607.500000 397.650000 649.500000 398.350000 ;
      RECT 557.500000 397.650000 599.500000 398.350000 ;
      RECT 507.500000 397.650000 549.500000 398.350000 ;
      RECT 457.500000 397.650000 499.500000 399.650000 ;
      RECT 407.500000 397.650000 449.500000 398.350000 ;
      RECT 357.500000 397.650000 399.500000 398.350000 ;
      RECT 307.500000 397.650000 349.500000 398.350000 ;
      RECT 257.500000 397.650000 299.500000 398.350000 ;
      RECT 207.500000 397.650000 249.500000 398.350000 ;
      RECT 157.500000 397.650000 199.500000 398.350000 ;
      RECT 107.500000 397.650000 149.500000 398.350000 ;
      RECT 57.500000 397.650000 99.500000 398.350000 ;
      RECT 15.500000 397.650000 49.500000 398.350000 ;
      RECT 1183.500000 396.350000 1183.980000 399.165000 ;
      RECT 1169.500000 396.350000 1170.500000 397.650000 ;
      RECT 1116.500000 396.350000 1149.500000 397.650000 ;
      RECT 1107.500000 396.350000 1108.500000 397.650000 ;
      RECT 1066.500000 396.350000 1099.500000 397.650000 ;
      RECT 1057.500000 396.350000 1058.500000 397.650000 ;
      RECT 1016.500000 396.350000 1049.500000 397.650000 ;
      RECT 1007.500000 396.350000 1008.500000 397.650000 ;
      RECT 966.500000 396.350000 999.500000 397.650000 ;
      RECT 957.500000 396.350000 958.500000 397.650000 ;
      RECT 916.500000 396.350000 949.500000 397.650000 ;
      RECT 907.500000 396.350000 908.500000 397.650000 ;
      RECT 866.500000 396.350000 899.500000 397.650000 ;
      RECT 857.500000 396.350000 858.500000 397.650000 ;
      RECT 816.500000 396.350000 849.500000 397.650000 ;
      RECT 807.500000 396.350000 808.500000 397.650000 ;
      RECT 766.500000 396.350000 799.500000 397.650000 ;
      RECT 757.500000 396.350000 758.500000 397.650000 ;
      RECT 716.500000 396.350000 749.500000 397.650000 ;
      RECT 707.500000 396.350000 708.500000 397.650000 ;
      RECT 666.500000 396.350000 699.500000 397.650000 ;
      RECT 657.500000 396.350000 658.500000 397.650000 ;
      RECT 616.500000 396.350000 649.500000 397.650000 ;
      RECT 607.500000 396.350000 608.500000 397.650000 ;
      RECT 566.500000 396.350000 599.500000 397.650000 ;
      RECT 557.500000 396.350000 558.500000 397.650000 ;
      RECT 516.500000 396.350000 549.500000 397.650000 ;
      RECT 507.500000 396.350000 508.500000 397.650000 ;
      RECT 466.500000 396.350000 499.500000 397.650000 ;
      RECT 457.500000 396.350000 458.500000 397.650000 ;
      RECT 416.500000 396.350000 449.500000 397.650000 ;
      RECT 407.500000 396.350000 408.500000 397.650000 ;
      RECT 366.500000 396.350000 399.500000 397.650000 ;
      RECT 357.500000 396.350000 358.500000 397.650000 ;
      RECT 316.500000 396.350000 349.500000 397.650000 ;
      RECT 307.500000 396.350000 308.500000 397.650000 ;
      RECT 266.500000 396.350000 299.500000 397.650000 ;
      RECT 257.500000 396.350000 258.500000 397.650000 ;
      RECT 216.500000 396.350000 249.500000 397.650000 ;
      RECT 207.500000 396.350000 208.500000 397.650000 ;
      RECT 166.500000 396.350000 199.500000 397.650000 ;
      RECT 157.500000 396.350000 158.500000 397.650000 ;
      RECT 116.500000 396.350000 149.500000 397.650000 ;
      RECT 107.500000 396.350000 108.500000 397.650000 ;
      RECT 66.500000 396.350000 99.500000 397.650000 ;
      RECT 57.500000 396.350000 58.500000 397.650000 ;
      RECT 29.500000 396.350000 49.500000 397.650000 ;
      RECT 15.500000 396.350000 16.500000 397.650000 ;
      RECT 2.020000 396.350000 2.500000 399.170000 ;
      RECT 2.020000 396.070000 16.500000 396.350000 ;
      RECT 1169.500000 396.065000 1183.980000 396.350000 ;
      RECT 1169.500000 395.650000 1186.000000 396.065000 ;
      RECT 1116.500000 395.650000 1156.500000 396.350000 ;
      RECT 1066.500000 395.650000 1108.500000 396.350000 ;
      RECT 1016.500000 395.650000 1058.500000 396.350000 ;
      RECT 966.500000 395.650000 1008.500000 396.350000 ;
      RECT 916.500000 395.650000 958.500000 396.350000 ;
      RECT 866.500000 395.650000 908.500000 396.350000 ;
      RECT 816.500000 395.650000 858.500000 396.350000 ;
      RECT 766.500000 395.650000 808.500000 396.350000 ;
      RECT 716.500000 395.650000 758.500000 396.350000 ;
      RECT 666.500000 395.650000 708.500000 396.350000 ;
      RECT 616.500000 395.650000 658.500000 396.350000 ;
      RECT 566.500000 395.650000 608.500000 396.350000 ;
      RECT 516.500000 395.650000 558.500000 396.350000 ;
      RECT 466.500000 395.650000 508.500000 396.350000 ;
      RECT 416.500000 395.650000 458.500000 396.350000 ;
      RECT 366.500000 395.650000 408.500000 396.350000 ;
      RECT 316.500000 395.650000 358.500000 396.350000 ;
      RECT 266.500000 395.650000 308.500000 396.350000 ;
      RECT 216.500000 395.650000 258.500000 396.350000 ;
      RECT 166.500000 395.650000 208.500000 396.350000 ;
      RECT 116.500000 395.650000 158.500000 396.350000 ;
      RECT 66.500000 395.650000 108.500000 396.350000 ;
      RECT 29.500000 395.650000 58.500000 396.350000 ;
      RECT 0.000000 395.650000 16.500000 396.070000 ;
      RECT 1169.500000 394.350000 1170.500000 395.650000 ;
      RECT 1116.500000 394.350000 1149.500000 395.650000 ;
      RECT 1107.500000 394.350000 1108.500000 395.650000 ;
      RECT 1066.500000 394.350000 1099.500000 395.650000 ;
      RECT 1057.500000 394.350000 1058.500000 395.650000 ;
      RECT 1016.500000 394.350000 1049.500000 395.650000 ;
      RECT 1007.500000 394.350000 1008.500000 395.650000 ;
      RECT 966.500000 394.350000 999.500000 395.650000 ;
      RECT 957.500000 394.350000 958.500000 395.650000 ;
      RECT 916.500000 394.350000 949.500000 395.650000 ;
      RECT 907.500000 394.350000 908.500000 395.650000 ;
      RECT 866.500000 394.350000 899.500000 395.650000 ;
      RECT 857.500000 394.350000 858.500000 395.650000 ;
      RECT 816.500000 394.350000 849.500000 395.650000 ;
      RECT 807.500000 394.350000 808.500000 395.650000 ;
      RECT 766.500000 394.350000 799.500000 395.650000 ;
      RECT 757.500000 394.350000 758.500000 395.650000 ;
      RECT 716.500000 394.350000 749.500000 395.650000 ;
      RECT 707.500000 394.350000 708.500000 395.650000 ;
      RECT 666.500000 394.350000 699.500000 395.650000 ;
      RECT 657.500000 394.350000 658.500000 395.650000 ;
      RECT 616.500000 394.350000 649.500000 395.650000 ;
      RECT 607.500000 394.350000 608.500000 395.650000 ;
      RECT 566.500000 394.350000 599.500000 395.650000 ;
      RECT 557.500000 394.350000 558.500000 395.650000 ;
      RECT 516.500000 394.350000 549.500000 395.650000 ;
      RECT 507.500000 394.350000 508.500000 395.650000 ;
      RECT 466.500000 394.350000 499.500000 395.650000 ;
      RECT 457.500000 394.350000 458.500000 395.650000 ;
      RECT 416.500000 394.350000 449.500000 395.650000 ;
      RECT 407.500000 394.350000 408.500000 395.650000 ;
      RECT 366.500000 394.350000 399.500000 395.650000 ;
      RECT 357.500000 394.350000 358.500000 395.650000 ;
      RECT 316.500000 394.350000 349.500000 395.650000 ;
      RECT 307.500000 394.350000 308.500000 395.650000 ;
      RECT 266.500000 394.350000 299.500000 395.650000 ;
      RECT 257.500000 394.350000 258.500000 395.650000 ;
      RECT 216.500000 394.350000 249.500000 395.650000 ;
      RECT 207.500000 394.350000 208.500000 395.650000 ;
      RECT 166.500000 394.350000 199.500000 395.650000 ;
      RECT 157.500000 394.350000 158.500000 395.650000 ;
      RECT 116.500000 394.350000 149.500000 395.650000 ;
      RECT 107.500000 394.350000 108.500000 395.650000 ;
      RECT 66.500000 394.350000 99.500000 395.650000 ;
      RECT 57.500000 394.350000 58.500000 395.650000 ;
      RECT 29.500000 394.350000 49.500000 395.650000 ;
      RECT 15.500000 394.350000 16.500000 395.650000 ;
      RECT 1157.500000 393.650000 1170.500000 394.350000 ;
      RECT 1107.500000 393.650000 1149.500000 394.350000 ;
      RECT 1057.500000 393.650000 1099.500000 394.350000 ;
      RECT 1007.500000 393.650000 1049.500000 394.350000 ;
      RECT 957.500000 393.650000 999.500000 394.350000 ;
      RECT 907.500000 393.650000 949.500000 394.350000 ;
      RECT 857.500000 393.650000 899.500000 394.350000 ;
      RECT 807.500000 393.650000 849.500000 394.350000 ;
      RECT 757.500000 393.650000 799.500000 394.350000 ;
      RECT 707.500000 393.650000 749.500000 394.350000 ;
      RECT 657.500000 393.650000 699.500000 394.350000 ;
      RECT 607.500000 393.650000 649.500000 394.350000 ;
      RECT 557.500000 393.650000 599.500000 394.350000 ;
      RECT 507.500000 393.650000 549.500000 394.350000 ;
      RECT 457.500000 393.650000 499.500000 394.350000 ;
      RECT 407.500000 393.650000 449.500000 394.350000 ;
      RECT 357.500000 393.650000 399.500000 394.350000 ;
      RECT 307.500000 393.650000 349.500000 394.350000 ;
      RECT 257.500000 393.650000 299.500000 394.350000 ;
      RECT 207.500000 393.650000 249.500000 394.350000 ;
      RECT 157.500000 393.650000 199.500000 394.350000 ;
      RECT 107.500000 393.650000 149.500000 394.350000 ;
      RECT 57.500000 393.650000 99.500000 394.350000 ;
      RECT 15.500000 393.650000 49.500000 394.350000 ;
      RECT 1183.500000 393.485000 1186.000000 395.650000 ;
      RECT 1183.500000 392.350000 1183.980000 393.485000 ;
      RECT 1169.500000 392.350000 1170.500000 393.650000 ;
      RECT 1116.500000 392.350000 1149.500000 393.650000 ;
      RECT 1107.500000 392.350000 1108.500000 393.650000 ;
      RECT 1066.500000 392.350000 1099.500000 393.650000 ;
      RECT 1057.500000 392.350000 1058.500000 393.650000 ;
      RECT 1016.500000 392.350000 1049.500000 393.650000 ;
      RECT 1007.500000 392.350000 1008.500000 393.650000 ;
      RECT 966.500000 392.350000 999.500000 393.650000 ;
      RECT 957.500000 392.350000 958.500000 393.650000 ;
      RECT 916.500000 392.350000 949.500000 393.650000 ;
      RECT 907.500000 392.350000 908.500000 393.650000 ;
      RECT 866.500000 392.350000 899.500000 393.650000 ;
      RECT 857.500000 392.350000 858.500000 393.650000 ;
      RECT 816.500000 392.350000 849.500000 393.650000 ;
      RECT 807.500000 392.350000 808.500000 393.650000 ;
      RECT 766.500000 392.350000 799.500000 393.650000 ;
      RECT 757.500000 392.350000 758.500000 393.650000 ;
      RECT 716.500000 392.350000 749.500000 393.650000 ;
      RECT 707.500000 392.350000 708.500000 393.650000 ;
      RECT 666.500000 392.350000 699.500000 393.650000 ;
      RECT 657.500000 392.350000 658.500000 393.650000 ;
      RECT 616.500000 392.350000 649.500000 393.650000 ;
      RECT 607.500000 392.350000 608.500000 393.650000 ;
      RECT 566.500000 392.350000 599.500000 393.650000 ;
      RECT 557.500000 392.350000 558.500000 393.650000 ;
      RECT 516.500000 392.350000 549.500000 393.650000 ;
      RECT 507.500000 392.350000 508.500000 393.650000 ;
      RECT 466.500000 392.350000 499.500000 393.650000 ;
      RECT 457.500000 392.350000 458.500000 393.650000 ;
      RECT 416.500000 392.350000 449.500000 393.650000 ;
      RECT 407.500000 392.350000 408.500000 393.650000 ;
      RECT 366.500000 392.350000 399.500000 393.650000 ;
      RECT 357.500000 392.350000 358.500000 393.650000 ;
      RECT 316.500000 392.350000 349.500000 393.650000 ;
      RECT 307.500000 392.350000 308.500000 393.650000 ;
      RECT 266.500000 392.350000 299.500000 393.650000 ;
      RECT 257.500000 392.350000 258.500000 393.650000 ;
      RECT 216.500000 392.350000 249.500000 393.650000 ;
      RECT 207.500000 392.350000 208.500000 393.650000 ;
      RECT 166.500000 392.350000 199.500000 393.650000 ;
      RECT 157.500000 392.350000 158.500000 393.650000 ;
      RECT 116.500000 392.350000 149.500000 393.650000 ;
      RECT 107.500000 392.350000 108.500000 393.650000 ;
      RECT 66.500000 392.350000 99.500000 393.650000 ;
      RECT 57.500000 392.350000 58.500000 393.650000 ;
      RECT 29.500000 392.350000 49.500000 393.650000 ;
      RECT 15.500000 392.350000 16.500000 393.650000 ;
      RECT 0.000000 392.350000 2.500000 395.650000 ;
      RECT 1169.500000 391.650000 1183.980000 392.350000 ;
      RECT 1116.500000 391.650000 1156.500000 392.350000 ;
      RECT 1066.500000 391.650000 1108.500000 392.350000 ;
      RECT 1016.500000 391.650000 1058.500000 392.350000 ;
      RECT 966.500000 391.650000 1008.500000 392.350000 ;
      RECT 916.500000 391.650000 958.500000 392.350000 ;
      RECT 866.500000 391.650000 908.500000 392.350000 ;
      RECT 816.500000 391.650000 858.500000 392.350000 ;
      RECT 766.500000 391.650000 808.500000 392.350000 ;
      RECT 716.500000 391.650000 758.500000 392.350000 ;
      RECT 666.500000 391.650000 708.500000 392.350000 ;
      RECT 616.500000 391.650000 658.500000 392.350000 ;
      RECT 566.500000 391.650000 608.500000 392.350000 ;
      RECT 516.500000 391.650000 558.500000 392.350000 ;
      RECT 466.500000 391.650000 508.500000 392.350000 ;
      RECT 416.500000 391.650000 458.500000 392.350000 ;
      RECT 366.500000 391.650000 408.500000 392.350000 ;
      RECT 316.500000 391.650000 358.500000 392.350000 ;
      RECT 266.500000 391.650000 308.500000 392.350000 ;
      RECT 216.500000 391.650000 258.500000 392.350000 ;
      RECT 166.500000 391.650000 208.500000 392.350000 ;
      RECT 116.500000 391.650000 158.500000 392.350000 ;
      RECT 66.500000 391.650000 108.500000 392.350000 ;
      RECT 29.500000 391.650000 58.500000 392.350000 ;
      RECT 0.000000 391.650000 16.500000 392.350000 ;
      RECT 1183.500000 390.385000 1183.980000 391.650000 ;
      RECT 1169.500000 390.350000 1170.500000 391.650000 ;
      RECT 1116.500000 390.350000 1149.500000 391.650000 ;
      RECT 1107.500000 390.350000 1108.500000 391.650000 ;
      RECT 1066.500000 390.350000 1099.500000 391.650000 ;
      RECT 1057.500000 390.350000 1058.500000 391.650000 ;
      RECT 1016.500000 390.350000 1049.500000 391.650000 ;
      RECT 1007.500000 390.350000 1008.500000 391.650000 ;
      RECT 966.500000 390.350000 999.500000 391.650000 ;
      RECT 957.500000 390.350000 958.500000 391.650000 ;
      RECT 916.500000 390.350000 949.500000 391.650000 ;
      RECT 907.500000 390.350000 908.500000 391.650000 ;
      RECT 866.500000 390.350000 899.500000 391.650000 ;
      RECT 857.500000 390.350000 858.500000 391.650000 ;
      RECT 816.500000 390.350000 849.500000 391.650000 ;
      RECT 807.500000 390.350000 808.500000 391.650000 ;
      RECT 766.500000 390.350000 799.500000 391.650000 ;
      RECT 757.500000 390.350000 758.500000 391.650000 ;
      RECT 716.500000 390.350000 749.500000 391.650000 ;
      RECT 707.500000 390.350000 708.500000 391.650000 ;
      RECT 666.500000 390.350000 699.500000 391.650000 ;
      RECT 657.500000 390.350000 658.500000 391.650000 ;
      RECT 616.500000 390.350000 649.500000 391.650000 ;
      RECT 607.500000 390.350000 608.500000 391.650000 ;
      RECT 566.500000 390.350000 599.500000 391.650000 ;
      RECT 557.500000 390.350000 558.500000 391.650000 ;
      RECT 516.500000 390.350000 549.500000 391.650000 ;
      RECT 507.500000 390.350000 508.500000 391.650000 ;
      RECT 466.500000 390.350000 499.500000 391.650000 ;
      RECT 457.500000 390.350000 458.500000 391.650000 ;
      RECT 416.500000 390.350000 449.500000 391.650000 ;
      RECT 407.500000 390.350000 408.500000 391.650000 ;
      RECT 366.500000 390.350000 399.500000 391.650000 ;
      RECT 357.500000 390.350000 358.500000 391.650000 ;
      RECT 316.500000 390.350000 349.500000 391.650000 ;
      RECT 307.500000 390.350000 308.500000 391.650000 ;
      RECT 266.500000 390.350000 299.500000 391.650000 ;
      RECT 257.500000 390.350000 258.500000 391.650000 ;
      RECT 216.500000 390.350000 249.500000 391.650000 ;
      RECT 207.500000 390.350000 208.500000 391.650000 ;
      RECT 166.500000 390.350000 199.500000 391.650000 ;
      RECT 157.500000 390.350000 158.500000 391.650000 ;
      RECT 116.500000 390.350000 149.500000 391.650000 ;
      RECT 107.500000 390.350000 108.500000 391.650000 ;
      RECT 66.500000 390.350000 99.500000 391.650000 ;
      RECT 57.500000 390.350000 58.500000 391.650000 ;
      RECT 29.500000 390.350000 49.500000 391.650000 ;
      RECT 15.500000 390.350000 16.500000 391.650000 ;
      RECT 1157.500000 389.650000 1170.500000 390.350000 ;
      RECT 1107.500000 389.650000 1149.500000 390.350000 ;
      RECT 1057.500000 389.650000 1099.500000 390.350000 ;
      RECT 1007.500000 389.650000 1049.500000 390.350000 ;
      RECT 957.500000 389.650000 999.500000 390.350000 ;
      RECT 907.500000 389.650000 949.500000 390.350000 ;
      RECT 857.500000 389.650000 899.500000 390.350000 ;
      RECT 807.500000 389.650000 849.500000 390.350000 ;
      RECT 757.500000 389.650000 799.500000 390.350000 ;
      RECT 707.500000 389.650000 749.500000 390.350000 ;
      RECT 657.500000 389.650000 699.500000 390.350000 ;
      RECT 607.500000 389.650000 649.500000 390.350000 ;
      RECT 557.500000 389.650000 599.500000 390.350000 ;
      RECT 507.500000 389.650000 549.500000 390.350000 ;
      RECT 457.500000 389.650000 499.500000 390.350000 ;
      RECT 407.500000 389.650000 449.500000 390.350000 ;
      RECT 357.500000 389.650000 399.500000 390.350000 ;
      RECT 307.500000 389.650000 349.500000 390.350000 ;
      RECT 257.500000 389.650000 299.500000 390.350000 ;
      RECT 207.500000 389.650000 249.500000 390.350000 ;
      RECT 157.500000 389.650000 199.500000 390.350000 ;
      RECT 107.500000 389.650000 149.500000 390.350000 ;
      RECT 57.500000 389.650000 99.500000 390.350000 ;
      RECT 15.500000 389.650000 49.500000 390.350000 ;
      RECT 1183.500000 389.525000 1186.000000 390.385000 ;
      RECT 0.000000 388.575000 2.500000 391.650000 ;
      RECT 1183.500000 388.350000 1183.980000 389.525000 ;
      RECT 1169.500000 388.350000 1170.500000 389.650000 ;
      RECT 1116.500000 388.350000 1149.500000 389.650000 ;
      RECT 1107.500000 388.350000 1108.500000 389.650000 ;
      RECT 1066.500000 388.350000 1099.500000 389.650000 ;
      RECT 1057.500000 388.350000 1058.500000 389.650000 ;
      RECT 1016.500000 388.350000 1049.500000 389.650000 ;
      RECT 1007.500000 388.350000 1008.500000 389.650000 ;
      RECT 966.500000 388.350000 999.500000 389.650000 ;
      RECT 957.500000 388.350000 958.500000 389.650000 ;
      RECT 916.500000 388.350000 949.500000 389.650000 ;
      RECT 907.500000 388.350000 908.500000 389.650000 ;
      RECT 866.500000 388.350000 899.500000 389.650000 ;
      RECT 857.500000 388.350000 858.500000 389.650000 ;
      RECT 816.500000 388.350000 849.500000 389.650000 ;
      RECT 807.500000 388.350000 808.500000 389.650000 ;
      RECT 766.500000 388.350000 799.500000 389.650000 ;
      RECT 757.500000 388.350000 758.500000 389.650000 ;
      RECT 716.500000 388.350000 749.500000 389.650000 ;
      RECT 707.500000 388.350000 708.500000 389.650000 ;
      RECT 666.500000 388.350000 699.500000 389.650000 ;
      RECT 657.500000 388.350000 658.500000 389.650000 ;
      RECT 616.500000 388.350000 649.500000 389.650000 ;
      RECT 607.500000 388.350000 608.500000 389.650000 ;
      RECT 566.500000 388.350000 599.500000 389.650000 ;
      RECT 557.500000 388.350000 558.500000 389.650000 ;
      RECT 516.500000 388.350000 549.500000 389.650000 ;
      RECT 507.500000 388.350000 508.500000 389.650000 ;
      RECT 466.500000 388.350000 499.500000 389.650000 ;
      RECT 457.500000 388.350000 458.500000 389.650000 ;
      RECT 416.500000 388.350000 449.500000 389.650000 ;
      RECT 407.500000 388.350000 408.500000 389.650000 ;
      RECT 366.500000 388.350000 399.500000 389.650000 ;
      RECT 357.500000 388.350000 358.500000 389.650000 ;
      RECT 316.500000 388.350000 349.500000 389.650000 ;
      RECT 307.500000 388.350000 308.500000 389.650000 ;
      RECT 266.500000 388.350000 299.500000 389.650000 ;
      RECT 257.500000 388.350000 258.500000 389.650000 ;
      RECT 216.500000 388.350000 249.500000 389.650000 ;
      RECT 207.500000 388.350000 208.500000 389.650000 ;
      RECT 166.500000 388.350000 199.500000 389.650000 ;
      RECT 157.500000 388.350000 158.500000 389.650000 ;
      RECT 116.500000 388.350000 149.500000 389.650000 ;
      RECT 107.500000 388.350000 108.500000 389.650000 ;
      RECT 66.500000 388.350000 99.500000 389.650000 ;
      RECT 57.500000 388.350000 58.500000 389.650000 ;
      RECT 29.500000 388.350000 49.500000 389.650000 ;
      RECT 15.500000 388.350000 16.500000 389.650000 ;
      RECT 2.020000 388.350000 2.500000 388.575000 ;
      RECT 1169.500000 387.650000 1183.980000 388.350000 ;
      RECT 1116.500000 387.650000 1156.500000 388.350000 ;
      RECT 1066.500000 387.650000 1108.500000 388.350000 ;
      RECT 1016.500000 387.650000 1058.500000 388.350000 ;
      RECT 966.500000 387.650000 1008.500000 388.350000 ;
      RECT 916.500000 387.650000 958.500000 388.350000 ;
      RECT 866.500000 387.650000 908.500000 388.350000 ;
      RECT 816.500000 387.650000 858.500000 388.350000 ;
      RECT 766.500000 387.650000 808.500000 388.350000 ;
      RECT 716.500000 387.650000 758.500000 388.350000 ;
      RECT 666.500000 387.650000 708.500000 388.350000 ;
      RECT 616.500000 387.650000 658.500000 388.350000 ;
      RECT 566.500000 387.650000 608.500000 388.350000 ;
      RECT 516.500000 387.650000 558.500000 388.350000 ;
      RECT 466.500000 387.650000 508.500000 388.350000 ;
      RECT 416.500000 387.650000 458.500000 388.350000 ;
      RECT 366.500000 387.650000 408.500000 388.350000 ;
      RECT 316.500000 387.650000 358.500000 388.350000 ;
      RECT 266.500000 387.650000 308.500000 388.350000 ;
      RECT 216.500000 387.650000 258.500000 388.350000 ;
      RECT 166.500000 387.650000 208.500000 388.350000 ;
      RECT 116.500000 387.650000 158.500000 388.350000 ;
      RECT 66.500000 387.650000 108.500000 388.350000 ;
      RECT 29.500000 387.650000 58.500000 388.350000 ;
      RECT 2.020000 387.650000 16.500000 388.350000 ;
      RECT 1183.500000 386.425000 1183.980000 387.650000 ;
      RECT 1169.500000 386.350000 1170.500000 387.650000 ;
      RECT 1116.500000 386.350000 1149.500000 387.650000 ;
      RECT 1107.500000 386.350000 1108.500000 387.650000 ;
      RECT 1066.500000 386.350000 1099.500000 387.650000 ;
      RECT 1057.500000 386.350000 1058.500000 387.650000 ;
      RECT 1016.500000 386.350000 1049.500000 387.650000 ;
      RECT 1007.500000 386.350000 1008.500000 387.650000 ;
      RECT 966.500000 386.350000 999.500000 387.650000 ;
      RECT 957.500000 386.350000 958.500000 387.650000 ;
      RECT 916.500000 386.350000 949.500000 387.650000 ;
      RECT 907.500000 386.350000 908.500000 387.650000 ;
      RECT 866.500000 386.350000 899.500000 387.650000 ;
      RECT 857.500000 386.350000 858.500000 387.650000 ;
      RECT 816.500000 386.350000 849.500000 387.650000 ;
      RECT 807.500000 386.350000 808.500000 387.650000 ;
      RECT 766.500000 386.350000 799.500000 387.650000 ;
      RECT 757.500000 386.350000 758.500000 387.650000 ;
      RECT 716.500000 386.350000 749.500000 387.650000 ;
      RECT 707.500000 386.350000 708.500000 387.650000 ;
      RECT 666.500000 386.350000 699.500000 387.650000 ;
      RECT 657.500000 386.350000 658.500000 387.650000 ;
      RECT 616.500000 386.350000 649.500000 387.650000 ;
      RECT 607.500000 386.350000 608.500000 387.650000 ;
      RECT 566.500000 386.350000 599.500000 387.650000 ;
      RECT 557.500000 386.350000 558.500000 387.650000 ;
      RECT 516.500000 386.350000 549.500000 387.650000 ;
      RECT 507.500000 386.350000 508.500000 387.650000 ;
      RECT 466.500000 386.350000 499.500000 387.650000 ;
      RECT 457.500000 386.350000 458.500000 387.650000 ;
      RECT 416.500000 386.350000 449.500000 387.650000 ;
      RECT 407.500000 386.350000 408.500000 387.650000 ;
      RECT 366.500000 386.350000 399.500000 387.650000 ;
      RECT 357.500000 386.350000 358.500000 387.650000 ;
      RECT 316.500000 386.350000 349.500000 387.650000 ;
      RECT 307.500000 386.350000 308.500000 387.650000 ;
      RECT 266.500000 386.350000 299.500000 387.650000 ;
      RECT 257.500000 386.350000 258.500000 387.650000 ;
      RECT 216.500000 386.350000 249.500000 387.650000 ;
      RECT 207.500000 386.350000 208.500000 387.650000 ;
      RECT 166.500000 386.350000 199.500000 387.650000 ;
      RECT 157.500000 386.350000 158.500000 387.650000 ;
      RECT 116.500000 386.350000 149.500000 387.650000 ;
      RECT 107.500000 386.350000 108.500000 387.650000 ;
      RECT 66.500000 386.350000 99.500000 387.650000 ;
      RECT 57.500000 386.350000 58.500000 387.650000 ;
      RECT 29.500000 386.350000 49.500000 387.650000 ;
      RECT 15.500000 386.350000 16.500000 387.650000 ;
      RECT 1157.500000 385.650000 1170.500000 386.350000 ;
      RECT 1107.500000 385.650000 1149.500000 386.350000 ;
      RECT 1057.500000 385.650000 1099.500000 386.350000 ;
      RECT 1007.500000 385.650000 1049.500000 386.350000 ;
      RECT 957.500000 385.650000 999.500000 386.350000 ;
      RECT 907.500000 385.650000 949.500000 386.350000 ;
      RECT 857.500000 385.650000 899.500000 386.350000 ;
      RECT 807.500000 385.650000 849.500000 386.350000 ;
      RECT 757.500000 385.650000 799.500000 386.350000 ;
      RECT 707.500000 385.650000 749.500000 386.350000 ;
      RECT 657.500000 385.650000 699.500000 386.350000 ;
      RECT 607.500000 385.650000 649.500000 386.350000 ;
      RECT 557.500000 385.650000 599.500000 386.350000 ;
      RECT 507.500000 385.650000 549.500000 386.350000 ;
      RECT 457.500000 385.650000 499.500000 386.350000 ;
      RECT 407.500000 385.650000 449.500000 386.350000 ;
      RECT 357.500000 385.650000 399.500000 386.350000 ;
      RECT 307.500000 385.650000 349.500000 386.350000 ;
      RECT 257.500000 385.650000 299.500000 386.350000 ;
      RECT 207.500000 385.650000 249.500000 386.350000 ;
      RECT 157.500000 385.650000 199.500000 386.350000 ;
      RECT 107.500000 385.650000 149.500000 386.350000 ;
      RECT 57.500000 385.650000 99.500000 386.350000 ;
      RECT 15.500000 385.650000 49.500000 386.350000 ;
      RECT 2.020000 385.475000 2.500000 387.650000 ;
      RECT 0.000000 384.615000 2.500000 385.475000 ;
      RECT 1183.500000 384.350000 1186.000000 386.425000 ;
      RECT 1169.500000 384.350000 1170.500000 385.650000 ;
      RECT 1116.500000 384.350000 1149.500000 385.650000 ;
      RECT 1107.500000 384.350000 1108.500000 385.650000 ;
      RECT 1066.500000 384.350000 1099.500000 385.650000 ;
      RECT 1057.500000 384.350000 1058.500000 385.650000 ;
      RECT 1016.500000 384.350000 1049.500000 385.650000 ;
      RECT 1007.500000 384.350000 1008.500000 385.650000 ;
      RECT 966.500000 384.350000 999.500000 385.650000 ;
      RECT 957.500000 384.350000 958.500000 385.650000 ;
      RECT 916.500000 384.350000 949.500000 385.650000 ;
      RECT 907.500000 384.350000 908.500000 385.650000 ;
      RECT 866.500000 384.350000 899.500000 385.650000 ;
      RECT 857.500000 384.350000 858.500000 385.650000 ;
      RECT 816.500000 384.350000 849.500000 385.650000 ;
      RECT 807.500000 384.350000 808.500000 385.650000 ;
      RECT 766.500000 384.350000 799.500000 385.650000 ;
      RECT 757.500000 384.350000 758.500000 385.650000 ;
      RECT 716.500000 384.350000 749.500000 385.650000 ;
      RECT 707.500000 384.350000 708.500000 385.650000 ;
      RECT 666.500000 384.350000 699.500000 385.650000 ;
      RECT 657.500000 384.350000 658.500000 385.650000 ;
      RECT 616.500000 384.350000 649.500000 385.650000 ;
      RECT 607.500000 384.350000 608.500000 385.650000 ;
      RECT 566.500000 384.350000 599.500000 385.650000 ;
      RECT 557.500000 384.350000 558.500000 385.650000 ;
      RECT 516.500000 384.350000 549.500000 385.650000 ;
      RECT 507.500000 384.350000 508.500000 385.650000 ;
      RECT 466.500000 384.350000 499.500000 385.650000 ;
      RECT 457.500000 384.350000 458.500000 385.650000 ;
      RECT 416.500000 384.350000 449.500000 385.650000 ;
      RECT 407.500000 384.350000 408.500000 385.650000 ;
      RECT 366.500000 384.350000 399.500000 385.650000 ;
      RECT 357.500000 384.350000 358.500000 385.650000 ;
      RECT 316.500000 384.350000 349.500000 385.650000 ;
      RECT 307.500000 384.350000 308.500000 385.650000 ;
      RECT 266.500000 384.350000 299.500000 385.650000 ;
      RECT 257.500000 384.350000 258.500000 385.650000 ;
      RECT 216.500000 384.350000 249.500000 385.650000 ;
      RECT 207.500000 384.350000 208.500000 385.650000 ;
      RECT 166.500000 384.350000 199.500000 385.650000 ;
      RECT 157.500000 384.350000 158.500000 385.650000 ;
      RECT 116.500000 384.350000 149.500000 385.650000 ;
      RECT 107.500000 384.350000 108.500000 385.650000 ;
      RECT 66.500000 384.350000 99.500000 385.650000 ;
      RECT 57.500000 384.350000 58.500000 385.650000 ;
      RECT 29.500000 384.350000 49.500000 385.650000 ;
      RECT 15.500000 384.350000 16.500000 385.650000 ;
      RECT 2.020000 384.350000 2.500000 384.615000 ;
      RECT 1169.500000 383.650000 1186.000000 384.350000 ;
      RECT 1116.500000 383.650000 1156.500000 384.350000 ;
      RECT 1066.500000 383.650000 1108.500000 384.350000 ;
      RECT 1016.500000 383.650000 1058.500000 384.350000 ;
      RECT 966.500000 383.650000 1008.500000 384.350000 ;
      RECT 916.500000 383.650000 958.500000 384.350000 ;
      RECT 866.500000 383.650000 908.500000 384.350000 ;
      RECT 816.500000 383.650000 858.500000 384.350000 ;
      RECT 766.500000 383.650000 808.500000 384.350000 ;
      RECT 716.500000 383.650000 758.500000 384.350000 ;
      RECT 666.500000 383.650000 708.500000 384.350000 ;
      RECT 616.500000 383.650000 658.500000 384.350000 ;
      RECT 566.500000 383.650000 608.500000 384.350000 ;
      RECT 516.500000 383.650000 558.500000 384.350000 ;
      RECT 466.500000 383.650000 508.500000 384.350000 ;
      RECT 416.500000 383.650000 458.500000 384.350000 ;
      RECT 366.500000 383.650000 408.500000 384.350000 ;
      RECT 316.500000 383.650000 358.500000 384.350000 ;
      RECT 266.500000 383.650000 308.500000 384.350000 ;
      RECT 216.500000 383.650000 258.500000 384.350000 ;
      RECT 166.500000 383.650000 208.500000 384.350000 ;
      RECT 116.500000 383.650000 158.500000 384.350000 ;
      RECT 66.500000 383.650000 108.500000 384.350000 ;
      RECT 29.500000 383.650000 58.500000 384.350000 ;
      RECT 2.020000 383.650000 16.500000 384.350000 ;
      RECT 1169.500000 382.350000 1170.500000 383.650000 ;
      RECT 1116.500000 382.350000 1149.500000 383.650000 ;
      RECT 1107.500000 382.350000 1108.500000 383.650000 ;
      RECT 1066.500000 382.350000 1099.500000 383.650000 ;
      RECT 1057.500000 382.350000 1058.500000 383.650000 ;
      RECT 1016.500000 382.350000 1049.500000 383.650000 ;
      RECT 1007.500000 382.350000 1008.500000 383.650000 ;
      RECT 966.500000 382.350000 999.500000 383.650000 ;
      RECT 957.500000 382.350000 958.500000 383.650000 ;
      RECT 916.500000 382.350000 949.500000 383.650000 ;
      RECT 907.500000 382.350000 908.500000 383.650000 ;
      RECT 866.500000 382.350000 899.500000 383.650000 ;
      RECT 857.500000 382.350000 858.500000 383.650000 ;
      RECT 816.500000 382.350000 849.500000 383.650000 ;
      RECT 807.500000 382.350000 808.500000 383.650000 ;
      RECT 766.500000 382.350000 799.500000 383.650000 ;
      RECT 757.500000 382.350000 758.500000 383.650000 ;
      RECT 716.500000 382.350000 749.500000 383.650000 ;
      RECT 707.500000 382.350000 708.500000 383.650000 ;
      RECT 666.500000 382.350000 699.500000 383.650000 ;
      RECT 657.500000 382.350000 658.500000 383.650000 ;
      RECT 616.500000 382.350000 649.500000 383.650000 ;
      RECT 607.500000 382.350000 608.500000 383.650000 ;
      RECT 566.500000 382.350000 599.500000 383.650000 ;
      RECT 557.500000 382.350000 558.500000 383.650000 ;
      RECT 516.500000 382.350000 549.500000 383.650000 ;
      RECT 507.500000 382.350000 508.500000 383.650000 ;
      RECT 466.500000 382.350000 499.500000 383.650000 ;
      RECT 457.500000 382.350000 458.500000 383.650000 ;
      RECT 416.500000 382.350000 449.500000 383.650000 ;
      RECT 407.500000 382.350000 408.500000 383.650000 ;
      RECT 366.500000 382.350000 399.500000 383.650000 ;
      RECT 357.500000 382.350000 358.500000 383.650000 ;
      RECT 316.500000 382.350000 349.500000 383.650000 ;
      RECT 307.500000 382.350000 308.500000 383.650000 ;
      RECT 266.500000 382.350000 299.500000 383.650000 ;
      RECT 257.500000 382.350000 258.500000 383.650000 ;
      RECT 216.500000 382.350000 249.500000 383.650000 ;
      RECT 207.500000 382.350000 208.500000 383.650000 ;
      RECT 166.500000 382.350000 199.500000 383.650000 ;
      RECT 157.500000 382.350000 158.500000 383.650000 ;
      RECT 116.500000 382.350000 149.500000 383.650000 ;
      RECT 107.500000 382.350000 108.500000 383.650000 ;
      RECT 66.500000 382.350000 99.500000 383.650000 ;
      RECT 57.500000 382.350000 58.500000 383.650000 ;
      RECT 29.500000 382.350000 49.500000 383.650000 ;
      RECT 15.500000 382.350000 16.500000 383.650000 ;
      RECT 1157.500000 381.650000 1170.500000 382.350000 ;
      RECT 1107.500000 381.650000 1149.500000 382.350000 ;
      RECT 1057.500000 381.650000 1099.500000 382.350000 ;
      RECT 1007.500000 381.650000 1049.500000 382.350000 ;
      RECT 957.500000 381.650000 999.500000 382.350000 ;
      RECT 907.500000 381.650000 949.500000 382.350000 ;
      RECT 857.500000 381.650000 899.500000 382.350000 ;
      RECT 807.500000 381.650000 849.500000 382.350000 ;
      RECT 757.500000 381.650000 799.500000 382.350000 ;
      RECT 707.500000 381.650000 749.500000 382.350000 ;
      RECT 657.500000 381.650000 699.500000 382.350000 ;
      RECT 607.500000 381.650000 649.500000 382.350000 ;
      RECT 557.500000 381.650000 599.500000 382.350000 ;
      RECT 507.500000 381.650000 549.500000 382.350000 ;
      RECT 457.500000 381.650000 499.500000 382.350000 ;
      RECT 407.500000 381.650000 449.500000 382.350000 ;
      RECT 357.500000 381.650000 399.500000 382.350000 ;
      RECT 307.500000 381.650000 349.500000 382.350000 ;
      RECT 257.500000 381.650000 299.500000 382.350000 ;
      RECT 207.500000 381.650000 249.500000 382.350000 ;
      RECT 157.500000 381.650000 199.500000 382.350000 ;
      RECT 107.500000 381.650000 149.500000 382.350000 ;
      RECT 57.500000 381.650000 99.500000 382.350000 ;
      RECT 15.500000 381.650000 49.500000 382.350000 ;
      RECT 2.020000 381.515000 2.500000 383.650000 ;
      RECT 1183.500000 380.350000 1186.000000 383.650000 ;
      RECT 1169.500000 380.350000 1170.500000 381.650000 ;
      RECT 1116.500000 380.350000 1149.500000 381.650000 ;
      RECT 1107.500000 380.350000 1108.500000 381.650000 ;
      RECT 1066.500000 380.350000 1099.500000 381.650000 ;
      RECT 1057.500000 380.350000 1058.500000 381.650000 ;
      RECT 1016.500000 380.350000 1049.500000 381.650000 ;
      RECT 1007.500000 380.350000 1008.500000 381.650000 ;
      RECT 966.500000 380.350000 999.500000 381.650000 ;
      RECT 957.500000 380.350000 958.500000 381.650000 ;
      RECT 916.500000 380.350000 949.500000 381.650000 ;
      RECT 907.500000 380.350000 908.500000 381.650000 ;
      RECT 866.500000 380.350000 899.500000 381.650000 ;
      RECT 857.500000 380.350000 858.500000 381.650000 ;
      RECT 816.500000 380.350000 849.500000 381.650000 ;
      RECT 807.500000 380.350000 808.500000 381.650000 ;
      RECT 766.500000 380.350000 799.500000 381.650000 ;
      RECT 757.500000 380.350000 758.500000 381.650000 ;
      RECT 716.500000 380.350000 749.500000 381.650000 ;
      RECT 707.500000 380.350000 708.500000 381.650000 ;
      RECT 666.500000 380.350000 699.500000 381.650000 ;
      RECT 657.500000 380.350000 658.500000 381.650000 ;
      RECT 616.500000 380.350000 649.500000 381.650000 ;
      RECT 607.500000 380.350000 608.500000 381.650000 ;
      RECT 566.500000 380.350000 599.500000 381.650000 ;
      RECT 557.500000 380.350000 558.500000 381.650000 ;
      RECT 516.500000 380.350000 549.500000 381.650000 ;
      RECT 507.500000 380.350000 508.500000 381.650000 ;
      RECT 466.500000 380.350000 499.500000 381.650000 ;
      RECT 457.500000 380.350000 458.500000 381.650000 ;
      RECT 416.500000 380.350000 449.500000 381.650000 ;
      RECT 407.500000 380.350000 408.500000 381.650000 ;
      RECT 366.500000 380.350000 399.500000 381.650000 ;
      RECT 357.500000 380.350000 358.500000 381.650000 ;
      RECT 316.500000 380.350000 349.500000 381.650000 ;
      RECT 307.500000 380.350000 308.500000 381.650000 ;
      RECT 266.500000 380.350000 299.500000 381.650000 ;
      RECT 257.500000 380.350000 258.500000 381.650000 ;
      RECT 216.500000 380.350000 249.500000 381.650000 ;
      RECT 207.500000 380.350000 208.500000 381.650000 ;
      RECT 166.500000 380.350000 199.500000 381.650000 ;
      RECT 157.500000 380.350000 158.500000 381.650000 ;
      RECT 116.500000 380.350000 149.500000 381.650000 ;
      RECT 107.500000 380.350000 108.500000 381.650000 ;
      RECT 66.500000 380.350000 99.500000 381.650000 ;
      RECT 57.500000 380.350000 58.500000 381.650000 ;
      RECT 29.500000 380.350000 49.500000 381.650000 ;
      RECT 15.500000 380.350000 16.500000 381.650000 ;
      RECT 0.000000 380.350000 2.500000 381.515000 ;
      RECT 1169.500000 379.650000 1186.000000 380.350000 ;
      RECT 1116.500000 379.650000 1156.500000 380.350000 ;
      RECT 1066.500000 379.650000 1108.500000 380.350000 ;
      RECT 1016.500000 379.650000 1058.500000 380.350000 ;
      RECT 966.500000 379.650000 1008.500000 380.350000 ;
      RECT 916.500000 379.650000 958.500000 380.350000 ;
      RECT 866.500000 379.650000 908.500000 380.350000 ;
      RECT 816.500000 379.650000 858.500000 380.350000 ;
      RECT 766.500000 379.650000 808.500000 380.350000 ;
      RECT 716.500000 379.650000 758.500000 380.350000 ;
      RECT 666.500000 379.650000 708.500000 380.350000 ;
      RECT 616.500000 379.650000 658.500000 380.350000 ;
      RECT 566.500000 379.650000 608.500000 380.350000 ;
      RECT 516.500000 379.650000 558.500000 380.350000 ;
      RECT 466.500000 379.650000 508.500000 380.350000 ;
      RECT 416.500000 379.650000 458.500000 380.350000 ;
      RECT 366.500000 379.650000 408.500000 380.350000 ;
      RECT 316.500000 379.650000 358.500000 380.350000 ;
      RECT 266.500000 379.650000 308.500000 380.350000 ;
      RECT 216.500000 379.650000 258.500000 380.350000 ;
      RECT 166.500000 379.650000 208.500000 380.350000 ;
      RECT 116.500000 379.650000 158.500000 380.350000 ;
      RECT 66.500000 379.650000 108.500000 380.350000 ;
      RECT 29.500000 379.650000 58.500000 380.350000 ;
      RECT 0.000000 379.650000 16.500000 380.350000 ;
      RECT 0.000000 378.935000 2.500000 379.650000 ;
      RECT 1183.500000 378.930000 1186.000000 379.650000 ;
      RECT 1169.500000 378.350000 1170.500000 379.650000 ;
      RECT 1116.500000 378.350000 1149.500000 379.650000 ;
      RECT 1107.500000 378.350000 1108.500000 379.650000 ;
      RECT 1066.500000 378.350000 1099.500000 379.650000 ;
      RECT 1057.500000 378.350000 1058.500000 379.650000 ;
      RECT 1016.500000 378.350000 1049.500000 379.650000 ;
      RECT 1007.500000 378.350000 1008.500000 379.650000 ;
      RECT 966.500000 378.350000 999.500000 379.650000 ;
      RECT 957.500000 378.350000 958.500000 379.650000 ;
      RECT 916.500000 378.350000 949.500000 379.650000 ;
      RECT 907.500000 378.350000 908.500000 379.650000 ;
      RECT 866.500000 378.350000 899.500000 379.650000 ;
      RECT 857.500000 378.350000 858.500000 379.650000 ;
      RECT 816.500000 378.350000 849.500000 379.650000 ;
      RECT 807.500000 378.350000 808.500000 379.650000 ;
      RECT 766.500000 378.350000 799.500000 379.650000 ;
      RECT 757.500000 378.350000 758.500000 379.650000 ;
      RECT 716.500000 378.350000 749.500000 379.650000 ;
      RECT 707.500000 378.350000 708.500000 379.650000 ;
      RECT 666.500000 378.350000 699.500000 379.650000 ;
      RECT 657.500000 378.350000 658.500000 379.650000 ;
      RECT 616.500000 378.350000 649.500000 379.650000 ;
      RECT 607.500000 378.350000 608.500000 379.650000 ;
      RECT 566.500000 378.350000 599.500000 379.650000 ;
      RECT 557.500000 378.350000 558.500000 379.650000 ;
      RECT 516.500000 378.350000 549.500000 379.650000 ;
      RECT 507.500000 378.350000 508.500000 379.650000 ;
      RECT 466.500000 378.350000 499.500000 379.650000 ;
      RECT 457.500000 378.350000 458.500000 379.650000 ;
      RECT 416.500000 378.350000 449.500000 379.650000 ;
      RECT 407.500000 378.350000 408.500000 379.650000 ;
      RECT 366.500000 378.350000 399.500000 379.650000 ;
      RECT 357.500000 378.350000 358.500000 379.650000 ;
      RECT 316.500000 378.350000 349.500000 379.650000 ;
      RECT 307.500000 378.350000 308.500000 379.650000 ;
      RECT 266.500000 378.350000 299.500000 379.650000 ;
      RECT 257.500000 378.350000 258.500000 379.650000 ;
      RECT 216.500000 378.350000 249.500000 379.650000 ;
      RECT 207.500000 378.350000 208.500000 379.650000 ;
      RECT 166.500000 378.350000 199.500000 379.650000 ;
      RECT 157.500000 378.350000 158.500000 379.650000 ;
      RECT 116.500000 378.350000 149.500000 379.650000 ;
      RECT 107.500000 378.350000 108.500000 379.650000 ;
      RECT 66.500000 378.350000 99.500000 379.650000 ;
      RECT 57.500000 378.350000 58.500000 379.650000 ;
      RECT 29.500000 378.350000 49.500000 379.650000 ;
      RECT 15.500000 378.350000 16.500000 379.650000 ;
      RECT 1157.500000 377.650000 1170.500000 378.350000 ;
      RECT 1107.500000 377.650000 1149.500000 378.350000 ;
      RECT 1057.500000 377.650000 1099.500000 378.350000 ;
      RECT 1007.500000 377.650000 1049.500000 378.350000 ;
      RECT 957.500000 377.650000 999.500000 378.350000 ;
      RECT 907.500000 377.650000 949.500000 378.350000 ;
      RECT 857.500000 377.650000 899.500000 378.350000 ;
      RECT 807.500000 377.650000 849.500000 378.350000 ;
      RECT 757.500000 377.650000 799.500000 378.350000 ;
      RECT 707.500000 377.650000 749.500000 378.350000 ;
      RECT 657.500000 377.650000 699.500000 378.350000 ;
      RECT 607.500000 377.650000 649.500000 378.350000 ;
      RECT 557.500000 377.650000 599.500000 378.350000 ;
      RECT 507.500000 377.650000 549.500000 378.350000 ;
      RECT 457.500000 377.650000 499.500000 378.350000 ;
      RECT 407.500000 377.650000 449.500000 378.350000 ;
      RECT 357.500000 377.650000 399.500000 378.350000 ;
      RECT 307.500000 377.650000 349.500000 378.350000 ;
      RECT 257.500000 377.650000 299.500000 378.350000 ;
      RECT 207.500000 377.650000 249.500000 378.350000 ;
      RECT 157.500000 377.650000 199.500000 378.350000 ;
      RECT 107.500000 377.650000 149.500000 378.350000 ;
      RECT 57.500000 377.650000 99.500000 378.350000 ;
      RECT 15.500000 377.650000 49.500000 378.350000 ;
      RECT 1183.500000 376.350000 1183.980000 378.930000 ;
      RECT 1169.500000 376.350000 1170.500000 377.650000 ;
      RECT 1116.500000 376.350000 1149.500000 377.650000 ;
      RECT 1107.500000 376.350000 1108.500000 377.650000 ;
      RECT 1066.500000 376.350000 1099.500000 377.650000 ;
      RECT 1057.500000 376.350000 1058.500000 377.650000 ;
      RECT 1016.500000 376.350000 1049.500000 377.650000 ;
      RECT 1007.500000 376.350000 1008.500000 377.650000 ;
      RECT 966.500000 376.350000 999.500000 377.650000 ;
      RECT 957.500000 376.350000 958.500000 377.650000 ;
      RECT 916.500000 376.350000 949.500000 377.650000 ;
      RECT 907.500000 376.350000 908.500000 377.650000 ;
      RECT 866.500000 376.350000 899.500000 377.650000 ;
      RECT 857.500000 376.350000 858.500000 377.650000 ;
      RECT 816.500000 376.350000 849.500000 377.650000 ;
      RECT 807.500000 376.350000 808.500000 377.650000 ;
      RECT 766.500000 376.350000 799.500000 377.650000 ;
      RECT 757.500000 376.350000 758.500000 377.650000 ;
      RECT 716.500000 376.350000 749.500000 377.650000 ;
      RECT 707.500000 376.350000 708.500000 377.650000 ;
      RECT 666.500000 376.350000 699.500000 377.650000 ;
      RECT 657.500000 376.350000 658.500000 377.650000 ;
      RECT 616.500000 376.350000 649.500000 377.650000 ;
      RECT 607.500000 376.350000 608.500000 377.650000 ;
      RECT 566.500000 376.350000 599.500000 377.650000 ;
      RECT 557.500000 376.350000 558.500000 377.650000 ;
      RECT 516.500000 376.350000 549.500000 377.650000 ;
      RECT 507.500000 376.350000 508.500000 377.650000 ;
      RECT 466.500000 376.350000 499.500000 377.650000 ;
      RECT 457.500000 376.350000 458.500000 377.650000 ;
      RECT 416.500000 376.350000 449.500000 377.650000 ;
      RECT 407.500000 376.350000 408.500000 377.650000 ;
      RECT 366.500000 376.350000 399.500000 377.650000 ;
      RECT 357.500000 376.350000 358.500000 377.650000 ;
      RECT 316.500000 376.350000 349.500000 377.650000 ;
      RECT 307.500000 376.350000 308.500000 377.650000 ;
      RECT 266.500000 376.350000 299.500000 377.650000 ;
      RECT 257.500000 376.350000 258.500000 377.650000 ;
      RECT 216.500000 376.350000 249.500000 377.650000 ;
      RECT 207.500000 376.350000 208.500000 377.650000 ;
      RECT 166.500000 376.350000 199.500000 377.650000 ;
      RECT 157.500000 376.350000 158.500000 377.650000 ;
      RECT 116.500000 376.350000 149.500000 377.650000 ;
      RECT 107.500000 376.350000 108.500000 377.650000 ;
      RECT 66.500000 376.350000 99.500000 377.650000 ;
      RECT 57.500000 376.350000 58.500000 377.650000 ;
      RECT 29.500000 376.350000 49.500000 377.650000 ;
      RECT 15.500000 376.350000 16.500000 377.650000 ;
      RECT 2.020000 376.350000 2.500000 378.935000 ;
      RECT 2.020000 375.835000 16.500000 376.350000 ;
      RECT 1169.500000 375.830000 1183.980000 376.350000 ;
      RECT 1169.500000 375.650000 1186.000000 375.830000 ;
      RECT 1116.500000 375.650000 1156.500000 376.350000 ;
      RECT 1066.500000 375.650000 1108.500000 376.350000 ;
      RECT 1016.500000 375.650000 1058.500000 376.350000 ;
      RECT 966.500000 375.650000 1008.500000 376.350000 ;
      RECT 916.500000 375.650000 958.500000 376.350000 ;
      RECT 866.500000 375.650000 908.500000 376.350000 ;
      RECT 816.500000 375.650000 858.500000 376.350000 ;
      RECT 766.500000 375.650000 808.500000 376.350000 ;
      RECT 716.500000 375.650000 758.500000 376.350000 ;
      RECT 666.500000 375.650000 708.500000 376.350000 ;
      RECT 616.500000 375.650000 658.500000 376.350000 ;
      RECT 566.500000 375.650000 608.500000 376.350000 ;
      RECT 516.500000 375.650000 558.500000 376.350000 ;
      RECT 466.500000 375.650000 508.500000 376.350000 ;
      RECT 416.500000 375.650000 458.500000 376.350000 ;
      RECT 366.500000 375.650000 408.500000 376.350000 ;
      RECT 316.500000 375.650000 358.500000 376.350000 ;
      RECT 266.500000 375.650000 308.500000 376.350000 ;
      RECT 216.500000 375.650000 258.500000 376.350000 ;
      RECT 166.500000 375.650000 208.500000 376.350000 ;
      RECT 116.500000 375.650000 158.500000 376.350000 ;
      RECT 66.500000 375.650000 108.500000 376.350000 ;
      RECT 29.500000 375.650000 58.500000 376.350000 ;
      RECT 0.000000 375.650000 16.500000 375.835000 ;
      RECT 1169.500000 374.350000 1170.500000 375.650000 ;
      RECT 1116.500000 374.350000 1149.500000 375.650000 ;
      RECT 1107.500000 374.350000 1108.500000 375.650000 ;
      RECT 1066.500000 374.350000 1099.500000 375.650000 ;
      RECT 1057.500000 374.350000 1058.500000 375.650000 ;
      RECT 1016.500000 374.350000 1049.500000 375.650000 ;
      RECT 1007.500000 374.350000 1008.500000 375.650000 ;
      RECT 966.500000 374.350000 999.500000 375.650000 ;
      RECT 957.500000 374.350000 958.500000 375.650000 ;
      RECT 916.500000 374.350000 949.500000 375.650000 ;
      RECT 907.500000 374.350000 908.500000 375.650000 ;
      RECT 866.500000 374.350000 899.500000 375.650000 ;
      RECT 857.500000 374.350000 858.500000 375.650000 ;
      RECT 816.500000 374.350000 849.500000 375.650000 ;
      RECT 807.500000 374.350000 808.500000 375.650000 ;
      RECT 766.500000 374.350000 799.500000 375.650000 ;
      RECT 757.500000 374.350000 758.500000 375.650000 ;
      RECT 716.500000 374.350000 749.500000 375.650000 ;
      RECT 707.500000 374.350000 708.500000 375.650000 ;
      RECT 666.500000 374.350000 699.500000 375.650000 ;
      RECT 657.500000 374.350000 658.500000 375.650000 ;
      RECT 616.500000 374.350000 649.500000 375.650000 ;
      RECT 607.500000 374.350000 608.500000 375.650000 ;
      RECT 566.500000 374.350000 599.500000 375.650000 ;
      RECT 557.500000 374.350000 558.500000 375.650000 ;
      RECT 516.500000 374.350000 549.500000 375.650000 ;
      RECT 507.500000 374.350000 508.500000 375.650000 ;
      RECT 466.500000 374.350000 499.500000 375.650000 ;
      RECT 457.500000 374.350000 458.500000 375.650000 ;
      RECT 416.500000 374.350000 449.500000 375.650000 ;
      RECT 407.500000 374.350000 408.500000 375.650000 ;
      RECT 366.500000 374.350000 399.500000 375.650000 ;
      RECT 357.500000 374.350000 358.500000 375.650000 ;
      RECT 316.500000 374.350000 349.500000 375.650000 ;
      RECT 307.500000 374.350000 308.500000 375.650000 ;
      RECT 266.500000 374.350000 299.500000 375.650000 ;
      RECT 257.500000 374.350000 258.500000 375.650000 ;
      RECT 216.500000 374.350000 249.500000 375.650000 ;
      RECT 207.500000 374.350000 208.500000 375.650000 ;
      RECT 166.500000 374.350000 199.500000 375.650000 ;
      RECT 157.500000 374.350000 158.500000 375.650000 ;
      RECT 116.500000 374.350000 149.500000 375.650000 ;
      RECT 107.500000 374.350000 108.500000 375.650000 ;
      RECT 66.500000 374.350000 99.500000 375.650000 ;
      RECT 57.500000 374.350000 58.500000 375.650000 ;
      RECT 29.500000 374.350000 49.500000 375.650000 ;
      RECT 15.500000 374.350000 16.500000 375.650000 ;
      RECT 1157.500000 373.650000 1170.500000 374.350000 ;
      RECT 1107.500000 373.650000 1149.500000 374.350000 ;
      RECT 1057.500000 373.650000 1099.500000 374.350000 ;
      RECT 1007.500000 373.650000 1049.500000 374.350000 ;
      RECT 957.500000 373.650000 999.500000 374.350000 ;
      RECT 907.500000 373.650000 949.500000 374.350000 ;
      RECT 857.500000 373.650000 899.500000 374.350000 ;
      RECT 807.500000 373.650000 849.500000 374.350000 ;
      RECT 757.500000 373.650000 799.500000 374.350000 ;
      RECT 707.500000 373.650000 749.500000 374.350000 ;
      RECT 657.500000 373.650000 699.500000 374.350000 ;
      RECT 607.500000 373.650000 649.500000 374.350000 ;
      RECT 557.500000 373.650000 599.500000 374.350000 ;
      RECT 507.500000 373.650000 549.500000 374.350000 ;
      RECT 457.500000 373.650000 499.500000 374.350000 ;
      RECT 407.500000 373.650000 449.500000 374.350000 ;
      RECT 357.500000 373.650000 399.500000 374.350000 ;
      RECT 307.500000 373.650000 349.500000 374.350000 ;
      RECT 257.500000 373.650000 299.500000 374.350000 ;
      RECT 207.500000 373.650000 249.500000 374.350000 ;
      RECT 157.500000 373.650000 199.500000 374.350000 ;
      RECT 107.500000 373.650000 149.500000 374.350000 ;
      RECT 57.500000 373.650000 99.500000 374.350000 ;
      RECT 15.500000 373.650000 49.500000 374.350000 ;
      RECT 1183.500000 372.350000 1186.000000 375.650000 ;
      RECT 1169.500000 372.350000 1170.500000 373.650000 ;
      RECT 1116.500000 372.350000 1149.500000 373.650000 ;
      RECT 1107.500000 372.350000 1108.500000 373.650000 ;
      RECT 1066.500000 372.350000 1099.500000 373.650000 ;
      RECT 1057.500000 372.350000 1058.500000 373.650000 ;
      RECT 1016.500000 372.350000 1049.500000 373.650000 ;
      RECT 1007.500000 372.350000 1008.500000 373.650000 ;
      RECT 966.500000 372.350000 999.500000 373.650000 ;
      RECT 957.500000 372.350000 958.500000 373.650000 ;
      RECT 916.500000 372.350000 949.500000 373.650000 ;
      RECT 907.500000 372.350000 908.500000 373.650000 ;
      RECT 866.500000 372.350000 899.500000 373.650000 ;
      RECT 857.500000 372.350000 858.500000 373.650000 ;
      RECT 816.500000 372.350000 849.500000 373.650000 ;
      RECT 807.500000 372.350000 808.500000 373.650000 ;
      RECT 766.500000 372.350000 799.500000 373.650000 ;
      RECT 757.500000 372.350000 758.500000 373.650000 ;
      RECT 716.500000 372.350000 749.500000 373.650000 ;
      RECT 707.500000 372.350000 708.500000 373.650000 ;
      RECT 666.500000 372.350000 699.500000 373.650000 ;
      RECT 657.500000 372.350000 658.500000 373.650000 ;
      RECT 616.500000 372.350000 649.500000 373.650000 ;
      RECT 607.500000 372.350000 608.500000 373.650000 ;
      RECT 566.500000 372.350000 599.500000 373.650000 ;
      RECT 557.500000 372.350000 558.500000 373.650000 ;
      RECT 516.500000 372.350000 549.500000 373.650000 ;
      RECT 507.500000 372.350000 508.500000 373.650000 ;
      RECT 466.500000 372.350000 499.500000 373.650000 ;
      RECT 457.500000 372.350000 458.500000 373.650000 ;
      RECT 416.500000 372.350000 449.500000 373.650000 ;
      RECT 407.500000 372.350000 408.500000 373.650000 ;
      RECT 366.500000 372.350000 399.500000 373.650000 ;
      RECT 357.500000 372.350000 358.500000 373.650000 ;
      RECT 316.500000 372.350000 349.500000 373.650000 ;
      RECT 307.500000 372.350000 308.500000 373.650000 ;
      RECT 266.500000 372.350000 299.500000 373.650000 ;
      RECT 257.500000 372.350000 258.500000 373.650000 ;
      RECT 216.500000 372.350000 249.500000 373.650000 ;
      RECT 207.500000 372.350000 208.500000 373.650000 ;
      RECT 166.500000 372.350000 199.500000 373.650000 ;
      RECT 157.500000 372.350000 158.500000 373.650000 ;
      RECT 116.500000 372.350000 149.500000 373.650000 ;
      RECT 107.500000 372.350000 108.500000 373.650000 ;
      RECT 66.500000 372.350000 99.500000 373.650000 ;
      RECT 57.500000 372.350000 58.500000 373.650000 ;
      RECT 29.500000 372.350000 49.500000 373.650000 ;
      RECT 15.500000 372.350000 16.500000 373.650000 ;
      RECT 0.000000 372.350000 2.500000 375.650000 ;
      RECT 1169.500000 371.650000 1186.000000 372.350000 ;
      RECT 1116.500000 371.650000 1156.500000 372.350000 ;
      RECT 1066.500000 371.650000 1108.500000 372.350000 ;
      RECT 1016.500000 371.650000 1058.500000 372.350000 ;
      RECT 966.500000 371.650000 1008.500000 372.350000 ;
      RECT 916.500000 371.650000 958.500000 372.350000 ;
      RECT 866.500000 371.650000 908.500000 372.350000 ;
      RECT 816.500000 371.650000 858.500000 372.350000 ;
      RECT 766.500000 371.650000 808.500000 372.350000 ;
      RECT 716.500000 371.650000 758.500000 372.350000 ;
      RECT 666.500000 371.650000 708.500000 372.350000 ;
      RECT 616.500000 371.650000 658.500000 372.350000 ;
      RECT 566.500000 371.650000 608.500000 372.350000 ;
      RECT 516.500000 371.650000 558.500000 372.350000 ;
      RECT 466.500000 371.650000 508.500000 372.350000 ;
      RECT 416.500000 371.650000 458.500000 372.350000 ;
      RECT 366.500000 371.650000 408.500000 372.350000 ;
      RECT 316.500000 371.650000 358.500000 372.350000 ;
      RECT 266.500000 371.650000 308.500000 372.350000 ;
      RECT 216.500000 371.650000 258.500000 372.350000 ;
      RECT 166.500000 371.650000 208.500000 372.350000 ;
      RECT 116.500000 371.650000 158.500000 372.350000 ;
      RECT 66.500000 371.650000 108.500000 372.350000 ;
      RECT 29.500000 371.650000 58.500000 372.350000 ;
      RECT 0.000000 371.650000 16.500000 372.350000 ;
      RECT 1169.500000 370.350000 1170.500000 371.650000 ;
      RECT 1116.500000 370.350000 1149.500000 371.650000 ;
      RECT 1107.500000 370.350000 1108.500000 371.650000 ;
      RECT 1066.500000 370.350000 1099.500000 371.650000 ;
      RECT 1057.500000 370.350000 1058.500000 371.650000 ;
      RECT 1016.500000 370.350000 1049.500000 371.650000 ;
      RECT 1007.500000 370.350000 1008.500000 371.650000 ;
      RECT 966.500000 370.350000 999.500000 371.650000 ;
      RECT 957.500000 370.350000 958.500000 371.650000 ;
      RECT 916.500000 370.350000 949.500000 371.650000 ;
      RECT 907.500000 370.350000 908.500000 371.650000 ;
      RECT 866.500000 370.350000 899.500000 371.650000 ;
      RECT 857.500000 370.350000 858.500000 371.650000 ;
      RECT 816.500000 370.350000 849.500000 371.650000 ;
      RECT 807.500000 370.350000 808.500000 371.650000 ;
      RECT 766.500000 370.350000 799.500000 371.650000 ;
      RECT 757.500000 370.350000 758.500000 371.650000 ;
      RECT 716.500000 370.350000 749.500000 371.650000 ;
      RECT 707.500000 370.350000 708.500000 371.650000 ;
      RECT 666.500000 370.350000 699.500000 371.650000 ;
      RECT 657.500000 370.350000 658.500000 371.650000 ;
      RECT 616.500000 370.350000 649.500000 371.650000 ;
      RECT 607.500000 370.350000 608.500000 371.650000 ;
      RECT 566.500000 370.350000 599.500000 371.650000 ;
      RECT 557.500000 370.350000 558.500000 371.650000 ;
      RECT 516.500000 370.350000 549.500000 371.650000 ;
      RECT 507.500000 370.350000 508.500000 371.650000 ;
      RECT 466.500000 370.350000 499.500000 371.650000 ;
      RECT 457.500000 370.350000 458.500000 371.650000 ;
      RECT 416.500000 370.350000 449.500000 371.650000 ;
      RECT 407.500000 370.350000 408.500000 371.650000 ;
      RECT 366.500000 370.350000 399.500000 371.650000 ;
      RECT 357.500000 370.350000 358.500000 371.650000 ;
      RECT 316.500000 370.350000 349.500000 371.650000 ;
      RECT 307.500000 370.350000 308.500000 371.650000 ;
      RECT 266.500000 370.350000 299.500000 371.650000 ;
      RECT 257.500000 370.350000 258.500000 371.650000 ;
      RECT 216.500000 370.350000 249.500000 371.650000 ;
      RECT 207.500000 370.350000 208.500000 371.650000 ;
      RECT 166.500000 370.350000 199.500000 371.650000 ;
      RECT 157.500000 370.350000 158.500000 371.650000 ;
      RECT 116.500000 370.350000 149.500000 371.650000 ;
      RECT 107.500000 370.350000 108.500000 371.650000 ;
      RECT 66.500000 370.350000 99.500000 371.650000 ;
      RECT 57.500000 370.350000 58.500000 371.650000 ;
      RECT 29.500000 370.350000 49.500000 371.650000 ;
      RECT 15.500000 370.350000 16.500000 371.650000 ;
      RECT 1157.500000 369.650000 1170.500000 370.350000 ;
      RECT 1107.500000 369.650000 1149.500000 370.350000 ;
      RECT 1057.500000 369.650000 1099.500000 370.350000 ;
      RECT 1007.500000 369.650000 1049.500000 370.350000 ;
      RECT 957.500000 369.650000 999.500000 370.350000 ;
      RECT 907.500000 369.650000 949.500000 370.350000 ;
      RECT 857.500000 369.650000 899.500000 370.350000 ;
      RECT 807.500000 369.650000 849.500000 370.350000 ;
      RECT 757.500000 369.650000 799.500000 370.350000 ;
      RECT 707.500000 369.650000 749.500000 370.350000 ;
      RECT 657.500000 369.650000 699.500000 370.350000 ;
      RECT 607.500000 369.650000 649.500000 370.350000 ;
      RECT 557.500000 369.650000 599.500000 370.350000 ;
      RECT 507.500000 369.650000 549.500000 370.350000 ;
      RECT 407.500000 369.650000 449.500000 370.350000 ;
      RECT 357.500000 369.650000 399.500000 370.350000 ;
      RECT 307.500000 369.650000 349.500000 370.350000 ;
      RECT 257.500000 369.650000 299.500000 370.350000 ;
      RECT 207.500000 369.650000 249.500000 370.350000 ;
      RECT 157.500000 369.650000 199.500000 370.350000 ;
      RECT 107.500000 369.650000 149.500000 370.350000 ;
      RECT 57.500000 369.650000 99.500000 370.350000 ;
      RECT 15.500000 369.650000 49.500000 370.350000 ;
      RECT 1183.500000 368.350000 1186.000000 371.650000 ;
      RECT 1169.500000 368.350000 1170.500000 369.650000 ;
      RECT 1116.500000 368.350000 1149.500000 369.650000 ;
      RECT 1107.500000 368.350000 1108.500000 369.650000 ;
      RECT 1066.500000 368.350000 1099.500000 369.650000 ;
      RECT 1057.500000 368.350000 1058.500000 369.650000 ;
      RECT 1016.500000 368.350000 1049.500000 369.650000 ;
      RECT 1007.500000 368.350000 1008.500000 369.650000 ;
      RECT 966.500000 368.350000 999.500000 369.650000 ;
      RECT 957.500000 368.350000 958.500000 369.650000 ;
      RECT 916.500000 368.350000 949.500000 369.650000 ;
      RECT 907.500000 368.350000 908.500000 369.650000 ;
      RECT 866.500000 368.350000 899.500000 369.650000 ;
      RECT 857.500000 368.350000 858.500000 369.650000 ;
      RECT 816.500000 368.350000 849.500000 369.650000 ;
      RECT 807.500000 368.350000 808.500000 369.650000 ;
      RECT 766.500000 368.350000 799.500000 369.650000 ;
      RECT 757.500000 368.350000 758.500000 369.650000 ;
      RECT 716.500000 368.350000 749.500000 369.650000 ;
      RECT 707.500000 368.350000 708.500000 369.650000 ;
      RECT 666.500000 368.350000 699.500000 369.650000 ;
      RECT 657.500000 368.350000 658.500000 369.650000 ;
      RECT 616.500000 368.350000 649.500000 369.650000 ;
      RECT 607.500000 368.350000 608.500000 369.650000 ;
      RECT 566.500000 368.350000 599.500000 369.650000 ;
      RECT 557.500000 368.350000 558.500000 369.650000 ;
      RECT 516.500000 368.350000 549.500000 369.650000 ;
      RECT 507.500000 368.350000 508.500000 369.650000 ;
      RECT 457.500000 368.350000 499.500000 370.350000 ;
      RECT 416.500000 368.350000 449.500000 369.650000 ;
      RECT 407.500000 368.350000 408.500000 369.650000 ;
      RECT 366.500000 368.350000 399.500000 369.650000 ;
      RECT 357.500000 368.350000 358.500000 369.650000 ;
      RECT 316.500000 368.350000 349.500000 369.650000 ;
      RECT 307.500000 368.350000 308.500000 369.650000 ;
      RECT 266.500000 368.350000 299.500000 369.650000 ;
      RECT 257.500000 368.350000 258.500000 369.650000 ;
      RECT 216.500000 368.350000 249.500000 369.650000 ;
      RECT 207.500000 368.350000 208.500000 369.650000 ;
      RECT 166.500000 368.350000 199.500000 369.650000 ;
      RECT 157.500000 368.350000 158.500000 369.650000 ;
      RECT 116.500000 368.350000 149.500000 369.650000 ;
      RECT 107.500000 368.350000 108.500000 369.650000 ;
      RECT 66.500000 368.350000 99.500000 369.650000 ;
      RECT 57.500000 368.350000 58.500000 369.650000 ;
      RECT 29.500000 368.350000 49.500000 369.650000 ;
      RECT 15.500000 368.350000 16.500000 369.650000 ;
      RECT 0.000000 368.350000 2.500000 371.650000 ;
      RECT 1169.500000 367.650000 1186.000000 368.350000 ;
      RECT 1116.500000 367.650000 1156.500000 368.350000 ;
      RECT 1066.500000 367.650000 1108.500000 368.350000 ;
      RECT 1016.500000 367.650000 1058.500000 368.350000 ;
      RECT 966.500000 367.650000 1008.500000 368.350000 ;
      RECT 916.500000 367.650000 958.500000 368.350000 ;
      RECT 866.500000 367.650000 908.500000 368.350000 ;
      RECT 816.500000 367.650000 858.500000 368.350000 ;
      RECT 766.500000 367.650000 808.500000 368.350000 ;
      RECT 716.500000 367.650000 758.500000 368.350000 ;
      RECT 666.500000 367.650000 708.500000 368.350000 ;
      RECT 616.500000 367.650000 658.500000 368.350000 ;
      RECT 566.500000 367.650000 608.500000 368.350000 ;
      RECT 516.500000 367.650000 558.500000 368.350000 ;
      RECT 416.500000 367.650000 508.500000 368.350000 ;
      RECT 366.500000 367.650000 408.500000 368.350000 ;
      RECT 316.500000 367.650000 358.500000 368.350000 ;
      RECT 266.500000 367.650000 308.500000 368.350000 ;
      RECT 216.500000 367.650000 258.500000 368.350000 ;
      RECT 166.500000 367.650000 208.500000 368.350000 ;
      RECT 116.500000 367.650000 158.500000 368.350000 ;
      RECT 66.500000 367.650000 108.500000 368.350000 ;
      RECT 29.500000 367.650000 58.500000 368.350000 ;
      RECT 0.000000 367.650000 16.500000 368.350000 ;
      RECT 1169.500000 366.350000 1170.500000 367.650000 ;
      RECT 1116.500000 366.350000 1149.500000 367.650000 ;
      RECT 1107.500000 366.350000 1108.500000 367.650000 ;
      RECT 1066.500000 366.350000 1099.500000 367.650000 ;
      RECT 1057.500000 366.350000 1058.500000 367.650000 ;
      RECT 1016.500000 366.350000 1049.500000 367.650000 ;
      RECT 1007.500000 366.350000 1008.500000 367.650000 ;
      RECT 966.500000 366.350000 999.500000 367.650000 ;
      RECT 957.500000 366.350000 958.500000 367.650000 ;
      RECT 916.500000 366.350000 949.500000 367.650000 ;
      RECT 907.500000 366.350000 908.500000 367.650000 ;
      RECT 866.500000 366.350000 899.500000 367.650000 ;
      RECT 857.500000 366.350000 858.500000 367.650000 ;
      RECT 816.500000 366.350000 849.500000 367.650000 ;
      RECT 807.500000 366.350000 808.500000 367.650000 ;
      RECT 766.500000 366.350000 799.500000 367.650000 ;
      RECT 757.500000 366.350000 758.500000 367.650000 ;
      RECT 716.500000 366.350000 749.500000 367.650000 ;
      RECT 707.500000 366.350000 708.500000 367.650000 ;
      RECT 666.500000 366.350000 699.500000 367.650000 ;
      RECT 657.500000 366.350000 658.500000 367.650000 ;
      RECT 616.500000 366.350000 649.500000 367.650000 ;
      RECT 607.500000 366.350000 608.500000 367.650000 ;
      RECT 566.500000 366.350000 599.500000 367.650000 ;
      RECT 557.500000 366.350000 558.500000 367.650000 ;
      RECT 516.500000 366.350000 549.500000 367.650000 ;
      RECT 507.500000 366.350000 508.500000 367.650000 ;
      RECT 416.500000 366.350000 499.500000 367.650000 ;
      RECT 407.500000 366.350000 408.500000 367.650000 ;
      RECT 366.500000 366.350000 399.500000 367.650000 ;
      RECT 357.500000 366.350000 358.500000 367.650000 ;
      RECT 316.500000 366.350000 349.500000 367.650000 ;
      RECT 307.500000 366.350000 308.500000 367.650000 ;
      RECT 266.500000 366.350000 299.500000 367.650000 ;
      RECT 257.500000 366.350000 258.500000 367.650000 ;
      RECT 216.500000 366.350000 249.500000 367.650000 ;
      RECT 207.500000 366.350000 208.500000 367.650000 ;
      RECT 166.500000 366.350000 199.500000 367.650000 ;
      RECT 157.500000 366.350000 158.500000 367.650000 ;
      RECT 116.500000 366.350000 149.500000 367.650000 ;
      RECT 107.500000 366.350000 108.500000 367.650000 ;
      RECT 66.500000 366.350000 99.500000 367.650000 ;
      RECT 57.500000 366.350000 58.500000 367.650000 ;
      RECT 29.500000 366.350000 49.500000 367.650000 ;
      RECT 15.500000 366.350000 16.500000 367.650000 ;
      RECT 1157.500000 365.650000 1170.500000 366.350000 ;
      RECT 1107.500000 365.650000 1149.500000 366.350000 ;
      RECT 1057.500000 365.650000 1099.500000 366.350000 ;
      RECT 1007.500000 365.650000 1049.500000 366.350000 ;
      RECT 957.500000 365.650000 999.500000 366.350000 ;
      RECT 907.500000 365.650000 949.500000 366.350000 ;
      RECT 857.500000 365.650000 899.500000 366.350000 ;
      RECT 807.500000 365.650000 849.500000 366.350000 ;
      RECT 757.500000 365.650000 799.500000 366.350000 ;
      RECT 707.500000 365.650000 749.500000 366.350000 ;
      RECT 657.500000 365.650000 699.500000 366.350000 ;
      RECT 607.500000 365.650000 649.500000 366.350000 ;
      RECT 557.500000 365.650000 599.500000 366.350000 ;
      RECT 507.500000 365.650000 549.500000 366.350000 ;
      RECT 407.500000 365.650000 499.500000 366.350000 ;
      RECT 357.500000 365.650000 399.500000 366.350000 ;
      RECT 307.500000 365.650000 349.500000 366.350000 ;
      RECT 257.500000 365.650000 299.500000 366.350000 ;
      RECT 207.500000 365.650000 249.500000 366.350000 ;
      RECT 157.500000 365.650000 199.500000 366.350000 ;
      RECT 107.500000 365.650000 149.500000 366.350000 ;
      RECT 57.500000 365.650000 99.500000 366.350000 ;
      RECT 15.500000 365.650000 49.500000 366.350000 ;
      RECT 1183.500000 364.350000 1186.000000 367.650000 ;
      RECT 1169.500000 364.350000 1170.500000 365.650000 ;
      RECT 1116.500000 364.350000 1149.500000 365.650000 ;
      RECT 1107.500000 364.350000 1108.500000 365.650000 ;
      RECT 1066.500000 364.350000 1099.500000 365.650000 ;
      RECT 1057.500000 364.350000 1058.500000 365.650000 ;
      RECT 1016.500000 364.350000 1049.500000 365.650000 ;
      RECT 1007.500000 364.350000 1008.500000 365.650000 ;
      RECT 966.500000 364.350000 999.500000 365.650000 ;
      RECT 957.500000 364.350000 958.500000 365.650000 ;
      RECT 916.500000 364.350000 949.500000 365.650000 ;
      RECT 907.500000 364.350000 908.500000 365.650000 ;
      RECT 866.500000 364.350000 899.500000 365.650000 ;
      RECT 857.500000 364.350000 858.500000 365.650000 ;
      RECT 816.500000 364.350000 849.500000 365.650000 ;
      RECT 807.500000 364.350000 808.500000 365.650000 ;
      RECT 766.500000 364.350000 799.500000 365.650000 ;
      RECT 757.500000 364.350000 758.500000 365.650000 ;
      RECT 716.500000 364.350000 749.500000 365.650000 ;
      RECT 707.500000 364.350000 708.500000 365.650000 ;
      RECT 666.500000 364.350000 699.500000 365.650000 ;
      RECT 657.500000 364.350000 658.500000 365.650000 ;
      RECT 616.500000 364.350000 649.500000 365.650000 ;
      RECT 607.500000 364.350000 608.500000 365.650000 ;
      RECT 566.500000 364.350000 599.500000 365.650000 ;
      RECT 557.500000 364.350000 558.500000 365.650000 ;
      RECT 516.500000 364.350000 549.500000 365.650000 ;
      RECT 507.500000 364.350000 508.500000 365.650000 ;
      RECT 416.500000 364.350000 499.500000 365.650000 ;
      RECT 407.500000 364.350000 408.500000 365.650000 ;
      RECT 366.500000 364.350000 399.500000 365.650000 ;
      RECT 357.500000 364.350000 358.500000 365.650000 ;
      RECT 316.500000 364.350000 349.500000 365.650000 ;
      RECT 307.500000 364.350000 308.500000 365.650000 ;
      RECT 266.500000 364.350000 299.500000 365.650000 ;
      RECT 257.500000 364.350000 258.500000 365.650000 ;
      RECT 216.500000 364.350000 249.500000 365.650000 ;
      RECT 207.500000 364.350000 208.500000 365.650000 ;
      RECT 166.500000 364.350000 199.500000 365.650000 ;
      RECT 157.500000 364.350000 158.500000 365.650000 ;
      RECT 116.500000 364.350000 149.500000 365.650000 ;
      RECT 107.500000 364.350000 108.500000 365.650000 ;
      RECT 66.500000 364.350000 99.500000 365.650000 ;
      RECT 57.500000 364.350000 58.500000 365.650000 ;
      RECT 29.500000 364.350000 49.500000 365.650000 ;
      RECT 15.500000 364.350000 16.500000 365.650000 ;
      RECT 0.000000 364.350000 2.500000 367.650000 ;
      RECT 1169.500000 363.650000 1186.000000 364.350000 ;
      RECT 1116.500000 363.650000 1156.500000 364.350000 ;
      RECT 1066.500000 363.650000 1108.500000 364.350000 ;
      RECT 1016.500000 363.650000 1058.500000 364.350000 ;
      RECT 966.500000 363.650000 1008.500000 364.350000 ;
      RECT 916.500000 363.650000 958.500000 364.350000 ;
      RECT 866.500000 363.650000 908.500000 364.350000 ;
      RECT 816.500000 363.650000 858.500000 364.350000 ;
      RECT 766.500000 363.650000 808.500000 364.350000 ;
      RECT 716.500000 363.650000 758.500000 364.350000 ;
      RECT 666.500000 363.650000 708.500000 364.350000 ;
      RECT 616.500000 363.650000 658.500000 364.350000 ;
      RECT 566.500000 363.650000 608.500000 364.350000 ;
      RECT 516.500000 363.650000 558.500000 364.350000 ;
      RECT 416.500000 363.650000 508.500000 364.350000 ;
      RECT 366.500000 363.650000 408.500000 364.350000 ;
      RECT 316.500000 363.650000 358.500000 364.350000 ;
      RECT 266.500000 363.650000 308.500000 364.350000 ;
      RECT 216.500000 363.650000 258.500000 364.350000 ;
      RECT 166.500000 363.650000 208.500000 364.350000 ;
      RECT 116.500000 363.650000 158.500000 364.350000 ;
      RECT 66.500000 363.650000 108.500000 364.350000 ;
      RECT 29.500000 363.650000 58.500000 364.350000 ;
      RECT 0.000000 363.650000 16.500000 364.350000 ;
      RECT 1169.500000 362.350000 1170.500000 363.650000 ;
      RECT 1116.500000 362.350000 1149.500000 363.650000 ;
      RECT 1107.500000 362.350000 1108.500000 363.650000 ;
      RECT 1066.500000 362.350000 1099.500000 363.650000 ;
      RECT 1057.500000 362.350000 1058.500000 363.650000 ;
      RECT 1016.500000 362.350000 1049.500000 363.650000 ;
      RECT 1007.500000 362.350000 1008.500000 363.650000 ;
      RECT 966.500000 362.350000 999.500000 363.650000 ;
      RECT 957.500000 362.350000 958.500000 363.650000 ;
      RECT 916.500000 362.350000 949.500000 363.650000 ;
      RECT 907.500000 362.350000 908.500000 363.650000 ;
      RECT 866.500000 362.350000 899.500000 363.650000 ;
      RECT 857.500000 362.350000 858.500000 363.650000 ;
      RECT 816.500000 362.350000 849.500000 363.650000 ;
      RECT 807.500000 362.350000 808.500000 363.650000 ;
      RECT 766.500000 362.350000 799.500000 363.650000 ;
      RECT 757.500000 362.350000 758.500000 363.650000 ;
      RECT 716.500000 362.350000 749.500000 363.650000 ;
      RECT 707.500000 362.350000 708.500000 363.650000 ;
      RECT 666.500000 362.350000 699.500000 363.650000 ;
      RECT 657.500000 362.350000 658.500000 363.650000 ;
      RECT 616.500000 362.350000 649.500000 363.650000 ;
      RECT 607.500000 362.350000 608.500000 363.650000 ;
      RECT 566.500000 362.350000 599.500000 363.650000 ;
      RECT 557.500000 362.350000 558.500000 363.650000 ;
      RECT 516.500000 362.350000 549.500000 363.650000 ;
      RECT 507.500000 362.350000 508.500000 363.650000 ;
      RECT 416.500000 362.350000 499.500000 363.650000 ;
      RECT 407.500000 362.350000 408.500000 363.650000 ;
      RECT 366.500000 362.350000 399.500000 363.650000 ;
      RECT 357.500000 362.350000 358.500000 363.650000 ;
      RECT 316.500000 362.350000 349.500000 363.650000 ;
      RECT 307.500000 362.350000 308.500000 363.650000 ;
      RECT 266.500000 362.350000 299.500000 363.650000 ;
      RECT 257.500000 362.350000 258.500000 363.650000 ;
      RECT 216.500000 362.350000 249.500000 363.650000 ;
      RECT 207.500000 362.350000 208.500000 363.650000 ;
      RECT 166.500000 362.350000 199.500000 363.650000 ;
      RECT 157.500000 362.350000 158.500000 363.650000 ;
      RECT 116.500000 362.350000 149.500000 363.650000 ;
      RECT 107.500000 362.350000 108.500000 363.650000 ;
      RECT 66.500000 362.350000 99.500000 363.650000 ;
      RECT 57.500000 362.350000 58.500000 363.650000 ;
      RECT 29.500000 362.350000 49.500000 363.650000 ;
      RECT 15.500000 362.350000 16.500000 363.650000 ;
      RECT 1157.500000 361.650000 1170.500000 362.350000 ;
      RECT 1107.500000 361.650000 1149.500000 362.350000 ;
      RECT 1057.500000 361.650000 1099.500000 362.350000 ;
      RECT 1007.500000 361.650000 1049.500000 362.350000 ;
      RECT 957.500000 361.650000 999.500000 362.350000 ;
      RECT 907.500000 361.650000 949.500000 362.350000 ;
      RECT 857.500000 361.650000 899.500000 362.350000 ;
      RECT 807.500000 361.650000 849.500000 362.350000 ;
      RECT 757.500000 361.650000 799.500000 362.350000 ;
      RECT 707.500000 361.650000 749.500000 362.350000 ;
      RECT 657.500000 361.650000 699.500000 362.350000 ;
      RECT 607.500000 361.650000 649.500000 362.350000 ;
      RECT 557.500000 361.650000 599.500000 362.350000 ;
      RECT 507.500000 361.650000 549.500000 362.350000 ;
      RECT 407.500000 361.650000 499.500000 362.350000 ;
      RECT 357.500000 361.650000 399.500000 362.350000 ;
      RECT 307.500000 361.650000 349.500000 362.350000 ;
      RECT 257.500000 361.650000 299.500000 362.350000 ;
      RECT 207.500000 361.650000 249.500000 362.350000 ;
      RECT 157.500000 361.650000 199.500000 362.350000 ;
      RECT 107.500000 361.650000 149.500000 362.350000 ;
      RECT 15.500000 361.650000 49.500000 362.350000 ;
      RECT 1183.500000 360.350000 1186.000000 363.650000 ;
      RECT 1169.500000 360.350000 1170.500000 361.650000 ;
      RECT 1116.500000 360.350000 1149.500000 361.650000 ;
      RECT 1107.500000 360.350000 1108.500000 361.650000 ;
      RECT 1066.500000 360.350000 1099.500000 361.650000 ;
      RECT 1057.500000 360.350000 1058.500000 361.650000 ;
      RECT 1016.500000 360.350000 1049.500000 361.650000 ;
      RECT 1007.500000 360.350000 1008.500000 361.650000 ;
      RECT 966.500000 360.350000 999.500000 361.650000 ;
      RECT 957.500000 360.350000 958.500000 361.650000 ;
      RECT 916.500000 360.350000 949.500000 361.650000 ;
      RECT 907.500000 360.350000 908.500000 361.650000 ;
      RECT 866.500000 360.350000 899.500000 361.650000 ;
      RECT 857.500000 360.350000 858.500000 361.650000 ;
      RECT 816.500000 360.350000 849.500000 361.650000 ;
      RECT 807.500000 360.350000 808.500000 361.650000 ;
      RECT 766.500000 360.350000 799.500000 361.650000 ;
      RECT 757.500000 360.350000 758.500000 361.650000 ;
      RECT 716.500000 360.350000 749.500000 361.650000 ;
      RECT 707.500000 360.350000 708.500000 361.650000 ;
      RECT 666.500000 360.350000 699.500000 361.650000 ;
      RECT 657.500000 360.350000 658.500000 361.650000 ;
      RECT 616.500000 360.350000 649.500000 361.650000 ;
      RECT 607.500000 360.350000 608.500000 361.650000 ;
      RECT 566.500000 360.350000 599.500000 361.650000 ;
      RECT 557.500000 360.350000 558.500000 361.650000 ;
      RECT 516.500000 360.350000 549.500000 361.650000 ;
      RECT 507.500000 360.350000 508.500000 361.650000 ;
      RECT 416.500000 360.350000 499.500000 361.650000 ;
      RECT 407.500000 360.350000 408.500000 361.650000 ;
      RECT 366.500000 360.350000 399.500000 361.650000 ;
      RECT 357.500000 360.350000 358.500000 361.650000 ;
      RECT 316.500000 360.350000 349.500000 361.650000 ;
      RECT 307.500000 360.350000 308.500000 361.650000 ;
      RECT 266.500000 360.350000 299.500000 361.650000 ;
      RECT 257.500000 360.350000 258.500000 361.650000 ;
      RECT 216.500000 360.350000 249.500000 361.650000 ;
      RECT 207.500000 360.350000 208.500000 361.650000 ;
      RECT 166.500000 360.350000 199.500000 361.650000 ;
      RECT 157.500000 360.350000 158.500000 361.650000 ;
      RECT 116.500000 360.350000 149.500000 361.650000 ;
      RECT 107.500000 360.350000 108.500000 361.650000 ;
      RECT 57.500000 360.350000 99.500000 362.350000 ;
      RECT 29.500000 360.350000 49.500000 361.650000 ;
      RECT 15.500000 360.350000 16.500000 361.650000 ;
      RECT 0.000000 360.350000 2.500000 363.650000 ;
      RECT 1169.500000 359.650000 1186.000000 360.350000 ;
      RECT 1116.500000 359.650000 1156.500000 360.350000 ;
      RECT 1066.500000 359.650000 1108.500000 360.350000 ;
      RECT 1016.500000 359.650000 1058.500000 360.350000 ;
      RECT 966.500000 359.650000 1008.500000 360.350000 ;
      RECT 916.500000 359.650000 958.500000 360.350000 ;
      RECT 866.500000 359.650000 908.500000 360.350000 ;
      RECT 816.500000 359.650000 858.500000 360.350000 ;
      RECT 766.500000 359.650000 808.500000 360.350000 ;
      RECT 716.500000 359.650000 758.500000 360.350000 ;
      RECT 666.500000 359.650000 708.500000 360.350000 ;
      RECT 616.500000 359.650000 658.500000 360.350000 ;
      RECT 566.500000 359.650000 608.500000 360.350000 ;
      RECT 516.500000 359.650000 558.500000 360.350000 ;
      RECT 416.500000 359.650000 508.500000 360.350000 ;
      RECT 366.500000 359.650000 408.500000 360.350000 ;
      RECT 316.500000 359.650000 358.500000 360.350000 ;
      RECT 266.500000 359.650000 308.500000 360.350000 ;
      RECT 216.500000 359.650000 258.500000 360.350000 ;
      RECT 166.500000 359.650000 208.500000 360.350000 ;
      RECT 116.500000 359.650000 158.500000 360.350000 ;
      RECT 29.500000 359.650000 108.500000 360.350000 ;
      RECT 0.000000 359.650000 16.500000 360.350000 ;
      RECT 1169.500000 358.350000 1170.500000 359.650000 ;
      RECT 1116.500000 358.350000 1149.500000 359.650000 ;
      RECT 1107.500000 358.350000 1108.500000 359.650000 ;
      RECT 1066.500000 358.350000 1099.500000 359.650000 ;
      RECT 1057.500000 358.350000 1058.500000 359.650000 ;
      RECT 1016.500000 358.350000 1049.500000 359.650000 ;
      RECT 1007.500000 358.350000 1008.500000 359.650000 ;
      RECT 966.500000 358.350000 999.500000 359.650000 ;
      RECT 957.500000 358.350000 958.500000 359.650000 ;
      RECT 916.500000 358.350000 949.500000 359.650000 ;
      RECT 907.500000 358.350000 908.500000 359.650000 ;
      RECT 866.500000 358.350000 899.500000 359.650000 ;
      RECT 857.500000 358.350000 858.500000 359.650000 ;
      RECT 816.500000 358.350000 849.500000 359.650000 ;
      RECT 807.500000 358.350000 808.500000 359.650000 ;
      RECT 766.500000 358.350000 799.500000 359.650000 ;
      RECT 757.500000 358.350000 758.500000 359.650000 ;
      RECT 716.500000 358.350000 749.500000 359.650000 ;
      RECT 707.500000 358.350000 708.500000 359.650000 ;
      RECT 666.500000 358.350000 699.500000 359.650000 ;
      RECT 657.500000 358.350000 658.500000 359.650000 ;
      RECT 616.500000 358.350000 649.500000 359.650000 ;
      RECT 607.500000 358.350000 608.500000 359.650000 ;
      RECT 566.500000 358.350000 599.500000 359.650000 ;
      RECT 557.500000 358.350000 558.500000 359.650000 ;
      RECT 516.500000 358.350000 549.500000 359.650000 ;
      RECT 507.500000 358.350000 508.500000 359.650000 ;
      RECT 416.500000 358.350000 499.500000 359.650000 ;
      RECT 407.500000 358.350000 408.500000 359.650000 ;
      RECT 366.500000 358.350000 399.500000 359.650000 ;
      RECT 357.500000 358.350000 358.500000 359.650000 ;
      RECT 316.500000 358.350000 349.500000 359.650000 ;
      RECT 307.500000 358.350000 308.500000 359.650000 ;
      RECT 266.500000 358.350000 299.500000 359.650000 ;
      RECT 257.500000 358.350000 258.500000 359.650000 ;
      RECT 216.500000 358.350000 249.500000 359.650000 ;
      RECT 207.500000 358.350000 208.500000 359.650000 ;
      RECT 166.500000 358.350000 199.500000 359.650000 ;
      RECT 157.500000 358.350000 158.500000 359.650000 ;
      RECT 116.500000 358.350000 149.500000 359.650000 ;
      RECT 107.500000 358.350000 108.500000 359.650000 ;
      RECT 29.500000 358.350000 99.500000 359.650000 ;
      RECT 15.500000 358.350000 16.500000 359.650000 ;
      RECT 1157.500000 357.650000 1170.500000 358.350000 ;
      RECT 1107.500000 357.650000 1149.500000 358.350000 ;
      RECT 1057.500000 357.650000 1099.500000 358.350000 ;
      RECT 1007.500000 357.650000 1049.500000 358.350000 ;
      RECT 957.500000 357.650000 999.500000 358.350000 ;
      RECT 907.500000 357.650000 949.500000 358.350000 ;
      RECT 857.500000 357.650000 899.500000 358.350000 ;
      RECT 807.500000 357.650000 849.500000 358.350000 ;
      RECT 757.500000 357.650000 799.500000 358.350000 ;
      RECT 707.500000 357.650000 749.500000 358.350000 ;
      RECT 657.500000 357.650000 699.500000 358.350000 ;
      RECT 607.500000 357.650000 649.500000 358.350000 ;
      RECT 557.500000 357.650000 599.500000 358.350000 ;
      RECT 507.500000 357.650000 549.500000 358.350000 ;
      RECT 407.500000 357.650000 499.500000 358.350000 ;
      RECT 357.500000 357.650000 399.500000 358.350000 ;
      RECT 307.500000 357.650000 349.500000 358.350000 ;
      RECT 257.500000 357.650000 299.500000 358.350000 ;
      RECT 207.500000 357.650000 249.500000 358.350000 ;
      RECT 157.500000 357.650000 199.500000 358.350000 ;
      RECT 107.500000 357.650000 149.500000 358.350000 ;
      RECT 15.500000 357.650000 99.500000 358.350000 ;
      RECT 1183.500000 356.350000 1186.000000 359.650000 ;
      RECT 1169.500000 356.350000 1170.500000 357.650000 ;
      RECT 1116.500000 356.350000 1149.500000 357.650000 ;
      RECT 1107.500000 356.350000 1108.500000 357.650000 ;
      RECT 1066.500000 356.350000 1099.500000 357.650000 ;
      RECT 1057.500000 356.350000 1058.500000 357.650000 ;
      RECT 1016.500000 356.350000 1049.500000 357.650000 ;
      RECT 1007.500000 356.350000 1008.500000 357.650000 ;
      RECT 966.500000 356.350000 999.500000 357.650000 ;
      RECT 957.500000 356.350000 958.500000 357.650000 ;
      RECT 916.500000 356.350000 949.500000 357.650000 ;
      RECT 907.500000 356.350000 908.500000 357.650000 ;
      RECT 866.500000 356.350000 899.500000 357.650000 ;
      RECT 857.500000 356.350000 858.500000 357.650000 ;
      RECT 816.500000 356.350000 849.500000 357.650000 ;
      RECT 807.500000 356.350000 808.500000 357.650000 ;
      RECT 766.500000 356.350000 799.500000 357.650000 ;
      RECT 757.500000 356.350000 758.500000 357.650000 ;
      RECT 716.500000 356.350000 749.500000 357.650000 ;
      RECT 707.500000 356.350000 708.500000 357.650000 ;
      RECT 666.500000 356.350000 699.500000 357.650000 ;
      RECT 657.500000 356.350000 658.500000 357.650000 ;
      RECT 616.500000 356.350000 649.500000 357.650000 ;
      RECT 607.500000 356.350000 608.500000 357.650000 ;
      RECT 566.500000 356.350000 599.500000 357.650000 ;
      RECT 557.500000 356.350000 558.500000 357.650000 ;
      RECT 516.500000 356.350000 549.500000 357.650000 ;
      RECT 507.500000 356.350000 508.500000 357.650000 ;
      RECT 416.500000 356.350000 499.500000 357.650000 ;
      RECT 407.500000 356.350000 408.500000 357.650000 ;
      RECT 366.500000 356.350000 399.500000 357.650000 ;
      RECT 357.500000 356.350000 358.500000 357.650000 ;
      RECT 316.500000 356.350000 349.500000 357.650000 ;
      RECT 307.500000 356.350000 308.500000 357.650000 ;
      RECT 266.500000 356.350000 299.500000 357.650000 ;
      RECT 257.500000 356.350000 258.500000 357.650000 ;
      RECT 216.500000 356.350000 249.500000 357.650000 ;
      RECT 207.500000 356.350000 208.500000 357.650000 ;
      RECT 166.500000 356.350000 199.500000 357.650000 ;
      RECT 157.500000 356.350000 158.500000 357.650000 ;
      RECT 116.500000 356.350000 149.500000 357.650000 ;
      RECT 107.500000 356.350000 108.500000 357.650000 ;
      RECT 29.500000 356.350000 99.500000 357.650000 ;
      RECT 15.500000 356.350000 16.500000 357.650000 ;
      RECT 0.000000 356.350000 2.500000 359.650000 ;
      RECT 1169.500000 355.650000 1186.000000 356.350000 ;
      RECT 1116.500000 355.650000 1156.500000 356.350000 ;
      RECT 1066.500000 355.650000 1108.500000 356.350000 ;
      RECT 1016.500000 355.650000 1058.500000 356.350000 ;
      RECT 966.500000 355.650000 1008.500000 356.350000 ;
      RECT 916.500000 355.650000 958.500000 356.350000 ;
      RECT 866.500000 355.650000 908.500000 356.350000 ;
      RECT 816.500000 355.650000 858.500000 356.350000 ;
      RECT 766.500000 355.650000 808.500000 356.350000 ;
      RECT 716.500000 355.650000 758.500000 356.350000 ;
      RECT 666.500000 355.650000 708.500000 356.350000 ;
      RECT 616.500000 355.650000 658.500000 356.350000 ;
      RECT 566.500000 355.650000 608.500000 356.350000 ;
      RECT 516.500000 355.650000 558.500000 356.350000 ;
      RECT 416.500000 355.650000 508.500000 356.350000 ;
      RECT 366.500000 355.650000 408.500000 356.350000 ;
      RECT 316.500000 355.650000 358.500000 356.350000 ;
      RECT 266.500000 355.650000 308.500000 356.350000 ;
      RECT 216.500000 355.650000 258.500000 356.350000 ;
      RECT 166.500000 355.650000 208.500000 356.350000 ;
      RECT 116.500000 355.650000 158.500000 356.350000 ;
      RECT 29.500000 355.650000 108.500000 356.350000 ;
      RECT 0.000000 355.650000 16.500000 356.350000 ;
      RECT 1169.500000 354.350000 1170.500000 355.650000 ;
      RECT 1116.500000 354.350000 1149.500000 355.650000 ;
      RECT 1107.500000 354.350000 1108.500000 355.650000 ;
      RECT 1066.500000 354.350000 1099.500000 355.650000 ;
      RECT 1057.500000 354.350000 1058.500000 355.650000 ;
      RECT 1016.500000 354.350000 1049.500000 355.650000 ;
      RECT 1007.500000 354.350000 1008.500000 355.650000 ;
      RECT 966.500000 354.350000 999.500000 355.650000 ;
      RECT 957.500000 354.350000 958.500000 355.650000 ;
      RECT 916.500000 354.350000 949.500000 355.650000 ;
      RECT 907.500000 354.350000 908.500000 355.650000 ;
      RECT 866.500000 354.350000 899.500000 355.650000 ;
      RECT 857.500000 354.350000 858.500000 355.650000 ;
      RECT 816.500000 354.350000 849.500000 355.650000 ;
      RECT 807.500000 354.350000 808.500000 355.650000 ;
      RECT 766.500000 354.350000 799.500000 355.650000 ;
      RECT 757.500000 354.350000 758.500000 355.650000 ;
      RECT 716.500000 354.350000 749.500000 355.650000 ;
      RECT 707.500000 354.350000 708.500000 355.650000 ;
      RECT 666.500000 354.350000 699.500000 355.650000 ;
      RECT 657.500000 354.350000 658.500000 355.650000 ;
      RECT 616.500000 354.350000 649.500000 355.650000 ;
      RECT 607.500000 354.350000 608.500000 355.650000 ;
      RECT 566.500000 354.350000 599.500000 355.650000 ;
      RECT 557.500000 354.350000 558.500000 355.650000 ;
      RECT 516.500000 354.350000 549.500000 355.650000 ;
      RECT 507.500000 354.350000 508.500000 355.650000 ;
      RECT 416.500000 354.350000 499.500000 355.650000 ;
      RECT 407.500000 354.350000 408.500000 355.650000 ;
      RECT 366.500000 354.350000 399.500000 355.650000 ;
      RECT 357.500000 354.350000 358.500000 355.650000 ;
      RECT 316.500000 354.350000 349.500000 355.650000 ;
      RECT 307.500000 354.350000 308.500000 355.650000 ;
      RECT 266.500000 354.350000 299.500000 355.650000 ;
      RECT 257.500000 354.350000 258.500000 355.650000 ;
      RECT 216.500000 354.350000 249.500000 355.650000 ;
      RECT 207.500000 354.350000 208.500000 355.650000 ;
      RECT 166.500000 354.350000 199.500000 355.650000 ;
      RECT 157.500000 354.350000 158.500000 355.650000 ;
      RECT 116.500000 354.350000 149.500000 355.650000 ;
      RECT 107.500000 354.350000 108.500000 355.650000 ;
      RECT 29.500000 354.350000 99.500000 355.650000 ;
      RECT 15.500000 354.350000 16.500000 355.650000 ;
      RECT 1157.500000 353.650000 1170.500000 354.350000 ;
      RECT 1107.500000 353.650000 1149.500000 354.350000 ;
      RECT 1057.500000 353.650000 1099.500000 354.350000 ;
      RECT 1007.500000 353.650000 1049.500000 354.350000 ;
      RECT 957.500000 353.650000 999.500000 354.350000 ;
      RECT 907.500000 353.650000 949.500000 354.350000 ;
      RECT 857.500000 353.650000 899.500000 354.350000 ;
      RECT 807.500000 353.650000 849.500000 354.350000 ;
      RECT 757.500000 353.650000 799.500000 354.350000 ;
      RECT 707.500000 353.650000 749.500000 354.350000 ;
      RECT 657.500000 353.650000 699.500000 354.350000 ;
      RECT 607.500000 353.650000 649.500000 354.350000 ;
      RECT 557.500000 353.650000 599.500000 354.350000 ;
      RECT 507.500000 353.650000 549.500000 354.350000 ;
      RECT 407.500000 353.650000 499.500000 354.350000 ;
      RECT 357.500000 353.650000 399.500000 354.350000 ;
      RECT 307.500000 353.650000 349.500000 354.350000 ;
      RECT 257.500000 353.650000 299.500000 354.350000 ;
      RECT 207.500000 353.650000 249.500000 354.350000 ;
      RECT 157.500000 353.650000 199.500000 354.350000 ;
      RECT 107.500000 353.650000 149.500000 354.350000 ;
      RECT 15.500000 353.650000 99.500000 354.350000 ;
      RECT 1183.500000 352.350000 1186.000000 355.650000 ;
      RECT 1169.500000 352.350000 1170.500000 353.650000 ;
      RECT 1116.500000 352.350000 1149.500000 353.650000 ;
      RECT 1107.500000 352.350000 1108.500000 353.650000 ;
      RECT 1066.500000 352.350000 1099.500000 353.650000 ;
      RECT 1057.500000 352.350000 1058.500000 353.650000 ;
      RECT 1016.500000 352.350000 1049.500000 353.650000 ;
      RECT 1007.500000 352.350000 1008.500000 353.650000 ;
      RECT 966.500000 352.350000 999.500000 353.650000 ;
      RECT 957.500000 352.350000 958.500000 353.650000 ;
      RECT 916.500000 352.350000 949.500000 353.650000 ;
      RECT 907.500000 352.350000 908.500000 353.650000 ;
      RECT 866.500000 352.350000 899.500000 353.650000 ;
      RECT 857.500000 352.350000 858.500000 353.650000 ;
      RECT 816.500000 352.350000 849.500000 353.650000 ;
      RECT 807.500000 352.350000 808.500000 353.650000 ;
      RECT 766.500000 352.350000 799.500000 353.650000 ;
      RECT 757.500000 352.350000 758.500000 353.650000 ;
      RECT 716.500000 352.350000 749.500000 353.650000 ;
      RECT 707.500000 352.350000 708.500000 353.650000 ;
      RECT 666.500000 352.350000 699.500000 353.650000 ;
      RECT 657.500000 352.350000 658.500000 353.650000 ;
      RECT 616.500000 352.350000 649.500000 353.650000 ;
      RECT 607.500000 352.350000 608.500000 353.650000 ;
      RECT 566.500000 352.350000 599.500000 353.650000 ;
      RECT 557.500000 352.350000 558.500000 353.650000 ;
      RECT 516.500000 352.350000 549.500000 353.650000 ;
      RECT 507.500000 352.350000 508.500000 353.650000 ;
      RECT 416.500000 352.350000 499.500000 353.650000 ;
      RECT 407.500000 352.350000 408.500000 353.650000 ;
      RECT 366.500000 352.350000 399.500000 353.650000 ;
      RECT 357.500000 352.350000 358.500000 353.650000 ;
      RECT 316.500000 352.350000 349.500000 353.650000 ;
      RECT 307.500000 352.350000 308.500000 353.650000 ;
      RECT 266.500000 352.350000 299.500000 353.650000 ;
      RECT 257.500000 352.350000 258.500000 353.650000 ;
      RECT 216.500000 352.350000 249.500000 353.650000 ;
      RECT 207.500000 352.350000 208.500000 353.650000 ;
      RECT 166.500000 352.350000 199.500000 353.650000 ;
      RECT 157.500000 352.350000 158.500000 353.650000 ;
      RECT 116.500000 352.350000 149.500000 353.650000 ;
      RECT 107.500000 352.350000 108.500000 353.650000 ;
      RECT 29.500000 352.350000 99.500000 353.650000 ;
      RECT 15.500000 352.350000 16.500000 353.650000 ;
      RECT 0.000000 352.350000 2.500000 355.650000 ;
      RECT 1169.500000 351.650000 1186.000000 352.350000 ;
      RECT 1116.500000 351.650000 1156.500000 352.350000 ;
      RECT 1066.500000 351.650000 1108.500000 352.350000 ;
      RECT 1016.500000 351.650000 1058.500000 352.350000 ;
      RECT 966.500000 351.650000 1008.500000 352.350000 ;
      RECT 916.500000 351.650000 958.500000 352.350000 ;
      RECT 866.500000 351.650000 908.500000 352.350000 ;
      RECT 816.500000 351.650000 858.500000 352.350000 ;
      RECT 766.500000 351.650000 808.500000 352.350000 ;
      RECT 716.500000 351.650000 758.500000 352.350000 ;
      RECT 666.500000 351.650000 708.500000 352.350000 ;
      RECT 616.500000 351.650000 658.500000 352.350000 ;
      RECT 566.500000 351.650000 608.500000 352.350000 ;
      RECT 516.500000 351.650000 558.500000 352.350000 ;
      RECT 416.500000 351.650000 508.500000 352.350000 ;
      RECT 366.500000 351.650000 408.500000 352.350000 ;
      RECT 316.500000 351.650000 358.500000 352.350000 ;
      RECT 266.500000 351.650000 308.500000 352.350000 ;
      RECT 216.500000 351.650000 258.500000 352.350000 ;
      RECT 166.500000 351.650000 208.500000 352.350000 ;
      RECT 116.500000 351.650000 158.500000 352.350000 ;
      RECT 29.500000 351.650000 108.500000 352.350000 ;
      RECT 0.000000 351.650000 16.500000 352.350000 ;
      RECT 1169.500000 350.350000 1170.500000 351.650000 ;
      RECT 1116.500000 350.350000 1149.500000 351.650000 ;
      RECT 1107.500000 350.350000 1108.500000 351.650000 ;
      RECT 1066.500000 350.350000 1099.500000 351.650000 ;
      RECT 1057.500000 350.350000 1058.500000 351.650000 ;
      RECT 1016.500000 350.350000 1049.500000 351.650000 ;
      RECT 1007.500000 350.350000 1008.500000 351.650000 ;
      RECT 966.500000 350.350000 999.500000 351.650000 ;
      RECT 957.500000 350.350000 958.500000 351.650000 ;
      RECT 916.500000 350.350000 949.500000 351.650000 ;
      RECT 907.500000 350.350000 908.500000 351.650000 ;
      RECT 866.500000 350.350000 899.500000 351.650000 ;
      RECT 857.500000 350.350000 858.500000 351.650000 ;
      RECT 816.500000 350.350000 849.500000 351.650000 ;
      RECT 807.500000 350.350000 808.500000 351.650000 ;
      RECT 766.500000 350.350000 799.500000 351.650000 ;
      RECT 757.500000 350.350000 758.500000 351.650000 ;
      RECT 716.500000 350.350000 749.500000 351.650000 ;
      RECT 707.500000 350.350000 708.500000 351.650000 ;
      RECT 666.500000 350.350000 699.500000 351.650000 ;
      RECT 657.500000 350.350000 658.500000 351.650000 ;
      RECT 616.500000 350.350000 649.500000 351.650000 ;
      RECT 607.500000 350.350000 608.500000 351.650000 ;
      RECT 566.500000 350.350000 599.500000 351.650000 ;
      RECT 557.500000 350.350000 558.500000 351.650000 ;
      RECT 516.500000 350.350000 549.500000 351.650000 ;
      RECT 507.500000 350.350000 508.500000 351.650000 ;
      RECT 416.500000 350.350000 499.500000 351.650000 ;
      RECT 407.500000 350.350000 408.500000 351.650000 ;
      RECT 366.500000 350.350000 399.500000 351.650000 ;
      RECT 357.500000 350.350000 358.500000 351.650000 ;
      RECT 316.500000 350.350000 349.500000 351.650000 ;
      RECT 307.500000 350.350000 308.500000 351.650000 ;
      RECT 266.500000 350.350000 299.500000 351.650000 ;
      RECT 257.500000 350.350000 258.500000 351.650000 ;
      RECT 216.500000 350.350000 249.500000 351.650000 ;
      RECT 207.500000 350.350000 208.500000 351.650000 ;
      RECT 166.500000 350.350000 199.500000 351.650000 ;
      RECT 157.500000 350.350000 158.500000 351.650000 ;
      RECT 116.500000 350.350000 149.500000 351.650000 ;
      RECT 107.500000 350.350000 108.500000 351.650000 ;
      RECT 29.500000 350.350000 99.500000 351.650000 ;
      RECT 15.500000 350.350000 16.500000 351.650000 ;
      RECT 1157.500000 349.650000 1170.500000 350.350000 ;
      RECT 1107.500000 349.650000 1149.500000 350.350000 ;
      RECT 1057.500000 349.650000 1099.500000 350.350000 ;
      RECT 1007.500000 349.650000 1049.500000 350.350000 ;
      RECT 957.500000 349.650000 999.500000 350.350000 ;
      RECT 907.500000 349.650000 949.500000 350.350000 ;
      RECT 857.500000 349.650000 899.500000 350.350000 ;
      RECT 807.500000 349.650000 849.500000 350.350000 ;
      RECT 757.500000 349.650000 799.500000 350.350000 ;
      RECT 707.500000 349.650000 749.500000 350.350000 ;
      RECT 657.500000 349.650000 699.500000 350.350000 ;
      RECT 607.500000 349.650000 649.500000 350.350000 ;
      RECT 557.500000 349.650000 599.500000 350.350000 ;
      RECT 507.500000 349.650000 549.500000 350.350000 ;
      RECT 407.500000 349.650000 499.500000 350.350000 ;
      RECT 357.500000 349.650000 399.500000 350.350000 ;
      RECT 307.500000 349.650000 349.500000 350.350000 ;
      RECT 257.500000 349.650000 299.500000 350.350000 ;
      RECT 207.500000 349.650000 249.500000 350.350000 ;
      RECT 157.500000 349.650000 199.500000 350.350000 ;
      RECT 107.500000 349.650000 149.500000 350.350000 ;
      RECT 15.500000 349.650000 99.500000 350.350000 ;
      RECT 1183.500000 348.350000 1186.000000 351.650000 ;
      RECT 1169.500000 348.350000 1170.500000 349.650000 ;
      RECT 1116.500000 348.350000 1149.500000 349.650000 ;
      RECT 1107.500000 348.350000 1108.500000 349.650000 ;
      RECT 1066.500000 348.350000 1099.500000 349.650000 ;
      RECT 1057.500000 348.350000 1058.500000 349.650000 ;
      RECT 1016.500000 348.350000 1049.500000 349.650000 ;
      RECT 1007.500000 348.350000 1008.500000 349.650000 ;
      RECT 966.500000 348.350000 999.500000 349.650000 ;
      RECT 957.500000 348.350000 958.500000 349.650000 ;
      RECT 916.500000 348.350000 949.500000 349.650000 ;
      RECT 907.500000 348.350000 908.500000 349.650000 ;
      RECT 866.500000 348.350000 899.500000 349.650000 ;
      RECT 857.500000 348.350000 858.500000 349.650000 ;
      RECT 816.500000 348.350000 849.500000 349.650000 ;
      RECT 807.500000 348.350000 808.500000 349.650000 ;
      RECT 766.500000 348.350000 799.500000 349.650000 ;
      RECT 757.500000 348.350000 758.500000 349.650000 ;
      RECT 716.500000 348.350000 749.500000 349.650000 ;
      RECT 707.500000 348.350000 708.500000 349.650000 ;
      RECT 666.500000 348.350000 699.500000 349.650000 ;
      RECT 657.500000 348.350000 658.500000 349.650000 ;
      RECT 616.500000 348.350000 649.500000 349.650000 ;
      RECT 607.500000 348.350000 608.500000 349.650000 ;
      RECT 566.500000 348.350000 599.500000 349.650000 ;
      RECT 557.500000 348.350000 558.500000 349.650000 ;
      RECT 516.500000 348.350000 549.500000 349.650000 ;
      RECT 507.500000 348.350000 508.500000 349.650000 ;
      RECT 466.500000 348.350000 499.500000 349.650000 ;
      RECT 407.500000 348.350000 408.500000 349.650000 ;
      RECT 366.500000 348.350000 399.500000 349.650000 ;
      RECT 357.500000 348.350000 358.500000 349.650000 ;
      RECT 316.500000 348.350000 349.500000 349.650000 ;
      RECT 307.500000 348.350000 308.500000 349.650000 ;
      RECT 266.500000 348.350000 299.500000 349.650000 ;
      RECT 257.500000 348.350000 258.500000 349.650000 ;
      RECT 216.500000 348.350000 249.500000 349.650000 ;
      RECT 207.500000 348.350000 208.500000 349.650000 ;
      RECT 166.500000 348.350000 199.500000 349.650000 ;
      RECT 157.500000 348.350000 158.500000 349.650000 ;
      RECT 116.500000 348.350000 149.500000 349.650000 ;
      RECT 107.500000 348.350000 108.500000 349.650000 ;
      RECT 66.500000 348.350000 99.500000 349.650000 ;
      RECT 15.500000 348.350000 16.500000 349.650000 ;
      RECT 0.000000 348.350000 2.500000 351.650000 ;
      RECT 1169.500000 347.650000 1186.000000 348.350000 ;
      RECT 1116.500000 347.650000 1156.500000 348.350000 ;
      RECT 1066.500000 347.650000 1108.500000 348.350000 ;
      RECT 1016.500000 347.650000 1058.500000 348.350000 ;
      RECT 966.500000 347.650000 1008.500000 348.350000 ;
      RECT 916.500000 347.650000 958.500000 348.350000 ;
      RECT 866.500000 347.650000 908.500000 348.350000 ;
      RECT 816.500000 347.650000 858.500000 348.350000 ;
      RECT 766.500000 347.650000 808.500000 348.350000 ;
      RECT 716.500000 347.650000 758.500000 348.350000 ;
      RECT 666.500000 347.650000 708.500000 348.350000 ;
      RECT 616.500000 347.650000 658.500000 348.350000 ;
      RECT 566.500000 347.650000 608.500000 348.350000 ;
      RECT 516.500000 347.650000 558.500000 348.350000 ;
      RECT 466.500000 347.650000 508.500000 348.350000 ;
      RECT 416.500000 347.650000 458.500000 349.650000 ;
      RECT 366.500000 347.650000 408.500000 348.350000 ;
      RECT 316.500000 347.650000 358.500000 348.350000 ;
      RECT 266.500000 347.650000 308.500000 348.350000 ;
      RECT 216.500000 347.650000 258.500000 348.350000 ;
      RECT 166.500000 347.650000 208.500000 348.350000 ;
      RECT 116.500000 347.650000 158.500000 348.350000 ;
      RECT 66.500000 347.650000 108.500000 348.350000 ;
      RECT 29.500000 347.650000 58.500000 349.650000 ;
      RECT 0.000000 347.650000 16.500000 348.350000 ;
      RECT 1169.500000 346.350000 1170.500000 347.650000 ;
      RECT 1116.500000 346.350000 1149.500000 347.650000 ;
      RECT 1107.500000 346.350000 1108.500000 347.650000 ;
      RECT 1066.500000 346.350000 1099.500000 347.650000 ;
      RECT 1057.500000 346.350000 1058.500000 347.650000 ;
      RECT 1016.500000 346.350000 1049.500000 347.650000 ;
      RECT 1007.500000 346.350000 1008.500000 347.650000 ;
      RECT 966.500000 346.350000 999.500000 347.650000 ;
      RECT 957.500000 346.350000 958.500000 347.650000 ;
      RECT 916.500000 346.350000 949.500000 347.650000 ;
      RECT 907.500000 346.350000 908.500000 347.650000 ;
      RECT 866.500000 346.350000 899.500000 347.650000 ;
      RECT 857.500000 346.350000 858.500000 347.650000 ;
      RECT 816.500000 346.350000 849.500000 347.650000 ;
      RECT 807.500000 346.350000 808.500000 347.650000 ;
      RECT 766.500000 346.350000 799.500000 347.650000 ;
      RECT 757.500000 346.350000 758.500000 347.650000 ;
      RECT 716.500000 346.350000 749.500000 347.650000 ;
      RECT 707.500000 346.350000 708.500000 347.650000 ;
      RECT 666.500000 346.350000 699.500000 347.650000 ;
      RECT 657.500000 346.350000 658.500000 347.650000 ;
      RECT 616.500000 346.350000 649.500000 347.650000 ;
      RECT 607.500000 346.350000 608.500000 347.650000 ;
      RECT 566.500000 346.350000 599.500000 347.650000 ;
      RECT 557.500000 346.350000 558.500000 347.650000 ;
      RECT 516.500000 346.350000 549.500000 347.650000 ;
      RECT 507.500000 346.350000 508.500000 347.650000 ;
      RECT 466.500000 346.350000 499.500000 347.650000 ;
      RECT 457.500000 346.350000 458.500000 347.650000 ;
      RECT 416.500000 346.350000 449.500000 347.650000 ;
      RECT 407.500000 346.350000 408.500000 347.650000 ;
      RECT 366.500000 346.350000 399.500000 347.650000 ;
      RECT 357.500000 346.350000 358.500000 347.650000 ;
      RECT 316.500000 346.350000 349.500000 347.650000 ;
      RECT 307.500000 346.350000 308.500000 347.650000 ;
      RECT 266.500000 346.350000 299.500000 347.650000 ;
      RECT 257.500000 346.350000 258.500000 347.650000 ;
      RECT 216.500000 346.350000 249.500000 347.650000 ;
      RECT 207.500000 346.350000 208.500000 347.650000 ;
      RECT 166.500000 346.350000 199.500000 347.650000 ;
      RECT 157.500000 346.350000 158.500000 347.650000 ;
      RECT 116.500000 346.350000 149.500000 347.650000 ;
      RECT 107.500000 346.350000 108.500000 347.650000 ;
      RECT 66.500000 346.350000 99.500000 347.650000 ;
      RECT 57.500000 346.350000 58.500000 347.650000 ;
      RECT 29.500000 346.350000 49.500000 347.650000 ;
      RECT 15.500000 346.350000 16.500000 347.650000 ;
      RECT 1157.500000 345.650000 1170.500000 346.350000 ;
      RECT 1107.500000 345.650000 1149.500000 346.350000 ;
      RECT 1057.500000 345.650000 1099.500000 346.350000 ;
      RECT 1007.500000 345.650000 1049.500000 346.350000 ;
      RECT 957.500000 345.650000 999.500000 346.350000 ;
      RECT 907.500000 345.650000 949.500000 346.350000 ;
      RECT 857.500000 345.650000 899.500000 346.350000 ;
      RECT 807.500000 345.650000 849.500000 346.350000 ;
      RECT 757.500000 345.650000 799.500000 346.350000 ;
      RECT 707.500000 345.650000 749.500000 346.350000 ;
      RECT 657.500000 345.650000 699.500000 346.350000 ;
      RECT 607.500000 345.650000 649.500000 346.350000 ;
      RECT 557.500000 345.650000 599.500000 346.350000 ;
      RECT 507.500000 345.650000 549.500000 346.350000 ;
      RECT 457.500000 345.650000 499.500000 346.350000 ;
      RECT 407.500000 345.650000 449.500000 346.350000 ;
      RECT 357.500000 345.650000 399.500000 346.350000 ;
      RECT 307.500000 345.650000 349.500000 346.350000 ;
      RECT 257.500000 345.650000 299.500000 346.350000 ;
      RECT 207.500000 345.650000 249.500000 346.350000 ;
      RECT 157.500000 345.650000 199.500000 346.350000 ;
      RECT 107.500000 345.650000 149.500000 346.350000 ;
      RECT 57.500000 345.650000 99.500000 346.350000 ;
      RECT 15.500000 345.650000 49.500000 346.350000 ;
      RECT 1183.500000 344.350000 1186.000000 347.650000 ;
      RECT 1169.500000 344.350000 1170.500000 345.650000 ;
      RECT 1116.500000 344.350000 1149.500000 345.650000 ;
      RECT 1107.500000 344.350000 1108.500000 345.650000 ;
      RECT 1066.500000 344.350000 1099.500000 345.650000 ;
      RECT 1057.500000 344.350000 1058.500000 345.650000 ;
      RECT 1016.500000 344.350000 1049.500000 345.650000 ;
      RECT 1007.500000 344.350000 1008.500000 345.650000 ;
      RECT 966.500000 344.350000 999.500000 345.650000 ;
      RECT 957.500000 344.350000 958.500000 345.650000 ;
      RECT 916.500000 344.350000 949.500000 345.650000 ;
      RECT 907.500000 344.350000 908.500000 345.650000 ;
      RECT 866.500000 344.350000 899.500000 345.650000 ;
      RECT 857.500000 344.350000 858.500000 345.650000 ;
      RECT 816.500000 344.350000 849.500000 345.650000 ;
      RECT 807.500000 344.350000 808.500000 345.650000 ;
      RECT 766.500000 344.350000 799.500000 345.650000 ;
      RECT 757.500000 344.350000 758.500000 345.650000 ;
      RECT 716.500000 344.350000 749.500000 345.650000 ;
      RECT 707.500000 344.350000 708.500000 345.650000 ;
      RECT 666.500000 344.350000 699.500000 345.650000 ;
      RECT 657.500000 344.350000 658.500000 345.650000 ;
      RECT 616.500000 344.350000 649.500000 345.650000 ;
      RECT 607.500000 344.350000 608.500000 345.650000 ;
      RECT 566.500000 344.350000 599.500000 345.650000 ;
      RECT 557.500000 344.350000 558.500000 345.650000 ;
      RECT 516.500000 344.350000 549.500000 345.650000 ;
      RECT 507.500000 344.350000 508.500000 345.650000 ;
      RECT 466.500000 344.350000 499.500000 345.650000 ;
      RECT 457.500000 344.350000 458.500000 345.650000 ;
      RECT 416.500000 344.350000 449.500000 345.650000 ;
      RECT 407.500000 344.350000 408.500000 345.650000 ;
      RECT 366.500000 344.350000 399.500000 345.650000 ;
      RECT 357.500000 344.350000 358.500000 345.650000 ;
      RECT 316.500000 344.350000 349.500000 345.650000 ;
      RECT 307.500000 344.350000 308.500000 345.650000 ;
      RECT 266.500000 344.350000 299.500000 345.650000 ;
      RECT 257.500000 344.350000 258.500000 345.650000 ;
      RECT 216.500000 344.350000 249.500000 345.650000 ;
      RECT 207.500000 344.350000 208.500000 345.650000 ;
      RECT 166.500000 344.350000 199.500000 345.650000 ;
      RECT 157.500000 344.350000 158.500000 345.650000 ;
      RECT 116.500000 344.350000 149.500000 345.650000 ;
      RECT 107.500000 344.350000 108.500000 345.650000 ;
      RECT 66.500000 344.350000 99.500000 345.650000 ;
      RECT 57.500000 344.350000 58.500000 345.650000 ;
      RECT 29.500000 344.350000 49.500000 345.650000 ;
      RECT 15.500000 344.350000 16.500000 345.650000 ;
      RECT 0.000000 344.350000 2.500000 347.650000 ;
      RECT 1169.500000 343.650000 1186.000000 344.350000 ;
      RECT 1116.500000 343.650000 1156.500000 344.350000 ;
      RECT 1066.500000 343.650000 1108.500000 344.350000 ;
      RECT 1016.500000 343.650000 1058.500000 344.350000 ;
      RECT 966.500000 343.650000 1008.500000 344.350000 ;
      RECT 916.500000 343.650000 958.500000 344.350000 ;
      RECT 866.500000 343.650000 908.500000 344.350000 ;
      RECT 816.500000 343.650000 858.500000 344.350000 ;
      RECT 766.500000 343.650000 808.500000 344.350000 ;
      RECT 716.500000 343.650000 758.500000 344.350000 ;
      RECT 666.500000 343.650000 708.500000 344.350000 ;
      RECT 616.500000 343.650000 658.500000 344.350000 ;
      RECT 566.500000 343.650000 608.500000 344.350000 ;
      RECT 516.500000 343.650000 558.500000 344.350000 ;
      RECT 466.500000 343.650000 508.500000 344.350000 ;
      RECT 416.500000 343.650000 458.500000 344.350000 ;
      RECT 366.500000 343.650000 408.500000 344.350000 ;
      RECT 316.500000 343.650000 358.500000 344.350000 ;
      RECT 266.500000 343.650000 308.500000 344.350000 ;
      RECT 216.500000 343.650000 258.500000 344.350000 ;
      RECT 166.500000 343.650000 208.500000 344.350000 ;
      RECT 116.500000 343.650000 158.500000 344.350000 ;
      RECT 66.500000 343.650000 108.500000 344.350000 ;
      RECT 29.500000 343.650000 58.500000 344.350000 ;
      RECT 0.000000 343.650000 16.500000 344.350000 ;
      RECT 1169.500000 342.350000 1170.500000 343.650000 ;
      RECT 1116.500000 342.350000 1149.500000 343.650000 ;
      RECT 1107.500000 342.350000 1108.500000 343.650000 ;
      RECT 1066.500000 342.350000 1099.500000 343.650000 ;
      RECT 1057.500000 342.350000 1058.500000 343.650000 ;
      RECT 1016.500000 342.350000 1049.500000 343.650000 ;
      RECT 1007.500000 342.350000 1008.500000 343.650000 ;
      RECT 966.500000 342.350000 999.500000 343.650000 ;
      RECT 957.500000 342.350000 958.500000 343.650000 ;
      RECT 916.500000 342.350000 949.500000 343.650000 ;
      RECT 907.500000 342.350000 908.500000 343.650000 ;
      RECT 866.500000 342.350000 899.500000 343.650000 ;
      RECT 857.500000 342.350000 858.500000 343.650000 ;
      RECT 816.500000 342.350000 849.500000 343.650000 ;
      RECT 807.500000 342.350000 808.500000 343.650000 ;
      RECT 766.500000 342.350000 799.500000 343.650000 ;
      RECT 757.500000 342.350000 758.500000 343.650000 ;
      RECT 716.500000 342.350000 749.500000 343.650000 ;
      RECT 707.500000 342.350000 708.500000 343.650000 ;
      RECT 666.500000 342.350000 699.500000 343.650000 ;
      RECT 657.500000 342.350000 658.500000 343.650000 ;
      RECT 616.500000 342.350000 649.500000 343.650000 ;
      RECT 607.500000 342.350000 608.500000 343.650000 ;
      RECT 566.500000 342.350000 599.500000 343.650000 ;
      RECT 557.500000 342.350000 558.500000 343.650000 ;
      RECT 516.500000 342.350000 549.500000 343.650000 ;
      RECT 507.500000 342.350000 508.500000 343.650000 ;
      RECT 466.500000 342.350000 499.500000 343.650000 ;
      RECT 457.500000 342.350000 458.500000 343.650000 ;
      RECT 416.500000 342.350000 449.500000 343.650000 ;
      RECT 407.500000 342.350000 408.500000 343.650000 ;
      RECT 366.500000 342.350000 399.500000 343.650000 ;
      RECT 357.500000 342.350000 358.500000 343.650000 ;
      RECT 316.500000 342.350000 349.500000 343.650000 ;
      RECT 307.500000 342.350000 308.500000 343.650000 ;
      RECT 266.500000 342.350000 299.500000 343.650000 ;
      RECT 257.500000 342.350000 258.500000 343.650000 ;
      RECT 216.500000 342.350000 249.500000 343.650000 ;
      RECT 207.500000 342.350000 208.500000 343.650000 ;
      RECT 166.500000 342.350000 199.500000 343.650000 ;
      RECT 157.500000 342.350000 158.500000 343.650000 ;
      RECT 116.500000 342.350000 149.500000 343.650000 ;
      RECT 107.500000 342.350000 108.500000 343.650000 ;
      RECT 66.500000 342.350000 99.500000 343.650000 ;
      RECT 57.500000 342.350000 58.500000 343.650000 ;
      RECT 29.500000 342.350000 49.500000 343.650000 ;
      RECT 15.500000 342.350000 16.500000 343.650000 ;
      RECT 1157.500000 341.650000 1170.500000 342.350000 ;
      RECT 1107.500000 341.650000 1149.500000 342.350000 ;
      RECT 1057.500000 341.650000 1099.500000 342.350000 ;
      RECT 1007.500000 341.650000 1049.500000 342.350000 ;
      RECT 957.500000 341.650000 999.500000 342.350000 ;
      RECT 907.500000 341.650000 949.500000 342.350000 ;
      RECT 857.500000 341.650000 899.500000 342.350000 ;
      RECT 807.500000 341.650000 849.500000 342.350000 ;
      RECT 757.500000 341.650000 799.500000 342.350000 ;
      RECT 707.500000 341.650000 749.500000 342.350000 ;
      RECT 657.500000 341.650000 699.500000 342.350000 ;
      RECT 607.500000 341.650000 649.500000 342.350000 ;
      RECT 557.500000 341.650000 599.500000 342.350000 ;
      RECT 507.500000 341.650000 549.500000 342.350000 ;
      RECT 457.500000 341.650000 499.500000 342.350000 ;
      RECT 407.500000 341.650000 449.500000 342.350000 ;
      RECT 357.500000 341.650000 399.500000 342.350000 ;
      RECT 307.500000 341.650000 349.500000 342.350000 ;
      RECT 257.500000 341.650000 299.500000 342.350000 ;
      RECT 207.500000 341.650000 249.500000 342.350000 ;
      RECT 157.500000 341.650000 199.500000 342.350000 ;
      RECT 107.500000 341.650000 149.500000 342.350000 ;
      RECT 57.500000 341.650000 99.500000 342.350000 ;
      RECT 15.500000 341.650000 49.500000 342.350000 ;
      RECT 1183.500000 340.350000 1186.000000 343.650000 ;
      RECT 1169.500000 340.350000 1170.500000 341.650000 ;
      RECT 1116.500000 340.350000 1149.500000 341.650000 ;
      RECT 1107.500000 340.350000 1108.500000 341.650000 ;
      RECT 1066.500000 340.350000 1099.500000 341.650000 ;
      RECT 1057.500000 340.350000 1058.500000 341.650000 ;
      RECT 1016.500000 340.350000 1049.500000 341.650000 ;
      RECT 1007.500000 340.350000 1008.500000 341.650000 ;
      RECT 966.500000 340.350000 999.500000 341.650000 ;
      RECT 957.500000 340.350000 958.500000 341.650000 ;
      RECT 916.500000 340.350000 949.500000 341.650000 ;
      RECT 907.500000 340.350000 908.500000 341.650000 ;
      RECT 866.500000 340.350000 899.500000 341.650000 ;
      RECT 857.500000 340.350000 858.500000 341.650000 ;
      RECT 816.500000 340.350000 849.500000 341.650000 ;
      RECT 807.500000 340.350000 808.500000 341.650000 ;
      RECT 766.500000 340.350000 799.500000 341.650000 ;
      RECT 757.500000 340.350000 758.500000 341.650000 ;
      RECT 716.500000 340.350000 749.500000 341.650000 ;
      RECT 707.500000 340.350000 708.500000 341.650000 ;
      RECT 666.500000 340.350000 699.500000 341.650000 ;
      RECT 657.500000 340.350000 658.500000 341.650000 ;
      RECT 616.500000 340.350000 649.500000 341.650000 ;
      RECT 607.500000 340.350000 608.500000 341.650000 ;
      RECT 566.500000 340.350000 599.500000 341.650000 ;
      RECT 557.500000 340.350000 558.500000 341.650000 ;
      RECT 516.500000 340.350000 549.500000 341.650000 ;
      RECT 507.500000 340.350000 508.500000 341.650000 ;
      RECT 466.500000 340.350000 499.500000 341.650000 ;
      RECT 457.500000 340.350000 458.500000 341.650000 ;
      RECT 416.500000 340.350000 449.500000 341.650000 ;
      RECT 407.500000 340.350000 408.500000 341.650000 ;
      RECT 366.500000 340.350000 399.500000 341.650000 ;
      RECT 357.500000 340.350000 358.500000 341.650000 ;
      RECT 316.500000 340.350000 349.500000 341.650000 ;
      RECT 307.500000 340.350000 308.500000 341.650000 ;
      RECT 266.500000 340.350000 299.500000 341.650000 ;
      RECT 257.500000 340.350000 258.500000 341.650000 ;
      RECT 216.500000 340.350000 249.500000 341.650000 ;
      RECT 207.500000 340.350000 208.500000 341.650000 ;
      RECT 166.500000 340.350000 199.500000 341.650000 ;
      RECT 157.500000 340.350000 158.500000 341.650000 ;
      RECT 116.500000 340.350000 149.500000 341.650000 ;
      RECT 107.500000 340.350000 108.500000 341.650000 ;
      RECT 66.500000 340.350000 99.500000 341.650000 ;
      RECT 57.500000 340.350000 58.500000 341.650000 ;
      RECT 29.500000 340.350000 49.500000 341.650000 ;
      RECT 15.500000 340.350000 16.500000 341.650000 ;
      RECT 0.000000 340.350000 2.500000 343.650000 ;
      RECT 1169.500000 339.650000 1186.000000 340.350000 ;
      RECT 1116.500000 339.650000 1156.500000 340.350000 ;
      RECT 1066.500000 339.650000 1108.500000 340.350000 ;
      RECT 1016.500000 339.650000 1058.500000 340.350000 ;
      RECT 966.500000 339.650000 1008.500000 340.350000 ;
      RECT 916.500000 339.650000 958.500000 340.350000 ;
      RECT 866.500000 339.650000 908.500000 340.350000 ;
      RECT 816.500000 339.650000 858.500000 340.350000 ;
      RECT 766.500000 339.650000 808.500000 340.350000 ;
      RECT 716.500000 339.650000 758.500000 340.350000 ;
      RECT 666.500000 339.650000 708.500000 340.350000 ;
      RECT 616.500000 339.650000 658.500000 340.350000 ;
      RECT 566.500000 339.650000 608.500000 340.350000 ;
      RECT 516.500000 339.650000 558.500000 340.350000 ;
      RECT 466.500000 339.650000 508.500000 340.350000 ;
      RECT 416.500000 339.650000 458.500000 340.350000 ;
      RECT 366.500000 339.650000 408.500000 340.350000 ;
      RECT 316.500000 339.650000 358.500000 340.350000 ;
      RECT 266.500000 339.650000 308.500000 340.350000 ;
      RECT 216.500000 339.650000 258.500000 340.350000 ;
      RECT 166.500000 339.650000 208.500000 340.350000 ;
      RECT 116.500000 339.650000 158.500000 340.350000 ;
      RECT 66.500000 339.650000 108.500000 340.350000 ;
      RECT 29.500000 339.650000 58.500000 340.350000 ;
      RECT 0.000000 339.650000 16.500000 340.350000 ;
      RECT 1169.500000 338.350000 1170.500000 339.650000 ;
      RECT 1116.500000 338.350000 1149.500000 339.650000 ;
      RECT 1107.500000 338.350000 1108.500000 339.650000 ;
      RECT 1066.500000 338.350000 1099.500000 339.650000 ;
      RECT 1057.500000 338.350000 1058.500000 339.650000 ;
      RECT 1016.500000 338.350000 1049.500000 339.650000 ;
      RECT 1007.500000 338.350000 1008.500000 339.650000 ;
      RECT 966.500000 338.350000 999.500000 339.650000 ;
      RECT 957.500000 338.350000 958.500000 339.650000 ;
      RECT 916.500000 338.350000 949.500000 339.650000 ;
      RECT 907.500000 338.350000 908.500000 339.650000 ;
      RECT 866.500000 338.350000 899.500000 339.650000 ;
      RECT 857.500000 338.350000 858.500000 339.650000 ;
      RECT 816.500000 338.350000 849.500000 339.650000 ;
      RECT 807.500000 338.350000 808.500000 339.650000 ;
      RECT 766.500000 338.350000 799.500000 339.650000 ;
      RECT 757.500000 338.350000 758.500000 339.650000 ;
      RECT 716.500000 338.350000 749.500000 339.650000 ;
      RECT 707.500000 338.350000 708.500000 339.650000 ;
      RECT 666.500000 338.350000 699.500000 339.650000 ;
      RECT 657.500000 338.350000 658.500000 339.650000 ;
      RECT 616.500000 338.350000 649.500000 339.650000 ;
      RECT 607.500000 338.350000 608.500000 339.650000 ;
      RECT 566.500000 338.350000 599.500000 339.650000 ;
      RECT 557.500000 338.350000 558.500000 339.650000 ;
      RECT 516.500000 338.350000 549.500000 339.650000 ;
      RECT 507.500000 338.350000 508.500000 339.650000 ;
      RECT 466.500000 338.350000 499.500000 339.650000 ;
      RECT 457.500000 338.350000 458.500000 339.650000 ;
      RECT 416.500000 338.350000 449.500000 339.650000 ;
      RECT 407.500000 338.350000 408.500000 339.650000 ;
      RECT 366.500000 338.350000 399.500000 339.650000 ;
      RECT 357.500000 338.350000 358.500000 339.650000 ;
      RECT 316.500000 338.350000 349.500000 339.650000 ;
      RECT 307.500000 338.350000 308.500000 339.650000 ;
      RECT 266.500000 338.350000 299.500000 339.650000 ;
      RECT 257.500000 338.350000 258.500000 339.650000 ;
      RECT 216.500000 338.350000 249.500000 339.650000 ;
      RECT 207.500000 338.350000 208.500000 339.650000 ;
      RECT 166.500000 338.350000 199.500000 339.650000 ;
      RECT 157.500000 338.350000 158.500000 339.650000 ;
      RECT 116.500000 338.350000 149.500000 339.650000 ;
      RECT 107.500000 338.350000 108.500000 339.650000 ;
      RECT 66.500000 338.350000 99.500000 339.650000 ;
      RECT 57.500000 338.350000 58.500000 339.650000 ;
      RECT 29.500000 338.350000 49.500000 339.650000 ;
      RECT 15.500000 338.350000 16.500000 339.650000 ;
      RECT 1157.500000 337.650000 1170.500000 338.350000 ;
      RECT 1107.500000 337.650000 1149.500000 338.350000 ;
      RECT 1057.500000 337.650000 1099.500000 338.350000 ;
      RECT 1007.500000 337.650000 1049.500000 338.350000 ;
      RECT 957.500000 337.650000 999.500000 338.350000 ;
      RECT 907.500000 337.650000 949.500000 338.350000 ;
      RECT 857.500000 337.650000 899.500000 338.350000 ;
      RECT 807.500000 337.650000 849.500000 338.350000 ;
      RECT 757.500000 337.650000 799.500000 338.350000 ;
      RECT 707.500000 337.650000 749.500000 338.350000 ;
      RECT 657.500000 337.650000 699.500000 338.350000 ;
      RECT 607.500000 337.650000 649.500000 338.350000 ;
      RECT 557.500000 337.650000 599.500000 338.350000 ;
      RECT 507.500000 337.650000 549.500000 338.350000 ;
      RECT 457.500000 337.650000 499.500000 338.350000 ;
      RECT 407.500000 337.650000 449.500000 338.350000 ;
      RECT 357.500000 337.650000 399.500000 338.350000 ;
      RECT 307.500000 337.650000 349.500000 338.350000 ;
      RECT 257.500000 337.650000 299.500000 338.350000 ;
      RECT 207.500000 337.650000 249.500000 338.350000 ;
      RECT 157.500000 337.650000 199.500000 338.350000 ;
      RECT 107.500000 337.650000 149.500000 338.350000 ;
      RECT 57.500000 337.650000 99.500000 338.350000 ;
      RECT 15.500000 337.650000 49.500000 338.350000 ;
      RECT 1183.500000 336.350000 1186.000000 339.650000 ;
      RECT 1169.500000 336.350000 1170.500000 337.650000 ;
      RECT 1116.500000 336.350000 1149.500000 337.650000 ;
      RECT 1107.500000 336.350000 1108.500000 337.650000 ;
      RECT 1066.500000 336.350000 1099.500000 337.650000 ;
      RECT 1057.500000 336.350000 1058.500000 337.650000 ;
      RECT 1016.500000 336.350000 1049.500000 337.650000 ;
      RECT 1007.500000 336.350000 1008.500000 337.650000 ;
      RECT 966.500000 336.350000 999.500000 337.650000 ;
      RECT 957.500000 336.350000 958.500000 337.650000 ;
      RECT 916.500000 336.350000 949.500000 337.650000 ;
      RECT 907.500000 336.350000 908.500000 337.650000 ;
      RECT 866.500000 336.350000 899.500000 337.650000 ;
      RECT 857.500000 336.350000 858.500000 337.650000 ;
      RECT 816.500000 336.350000 849.500000 337.650000 ;
      RECT 807.500000 336.350000 808.500000 337.650000 ;
      RECT 766.500000 336.350000 799.500000 337.650000 ;
      RECT 757.500000 336.350000 758.500000 337.650000 ;
      RECT 716.500000 336.350000 749.500000 337.650000 ;
      RECT 707.500000 336.350000 708.500000 337.650000 ;
      RECT 666.500000 336.350000 699.500000 337.650000 ;
      RECT 657.500000 336.350000 658.500000 337.650000 ;
      RECT 616.500000 336.350000 649.500000 337.650000 ;
      RECT 607.500000 336.350000 608.500000 337.650000 ;
      RECT 566.500000 336.350000 599.500000 337.650000 ;
      RECT 557.500000 336.350000 558.500000 337.650000 ;
      RECT 516.500000 336.350000 549.500000 337.650000 ;
      RECT 507.500000 336.350000 508.500000 337.650000 ;
      RECT 466.500000 336.350000 499.500000 337.650000 ;
      RECT 457.500000 336.350000 458.500000 337.650000 ;
      RECT 416.500000 336.350000 449.500000 337.650000 ;
      RECT 407.500000 336.350000 408.500000 337.650000 ;
      RECT 366.500000 336.350000 399.500000 337.650000 ;
      RECT 357.500000 336.350000 358.500000 337.650000 ;
      RECT 316.500000 336.350000 349.500000 337.650000 ;
      RECT 307.500000 336.350000 308.500000 337.650000 ;
      RECT 266.500000 336.350000 299.500000 337.650000 ;
      RECT 257.500000 336.350000 258.500000 337.650000 ;
      RECT 216.500000 336.350000 249.500000 337.650000 ;
      RECT 207.500000 336.350000 208.500000 337.650000 ;
      RECT 166.500000 336.350000 199.500000 337.650000 ;
      RECT 157.500000 336.350000 158.500000 337.650000 ;
      RECT 116.500000 336.350000 149.500000 337.650000 ;
      RECT 107.500000 336.350000 108.500000 337.650000 ;
      RECT 66.500000 336.350000 99.500000 337.650000 ;
      RECT 57.500000 336.350000 58.500000 337.650000 ;
      RECT 29.500000 336.350000 49.500000 337.650000 ;
      RECT 15.500000 336.350000 16.500000 337.650000 ;
      RECT 0.000000 336.350000 2.500000 339.650000 ;
      RECT 1169.500000 335.650000 1186.000000 336.350000 ;
      RECT 1116.500000 335.650000 1156.500000 336.350000 ;
      RECT 1066.500000 335.650000 1108.500000 336.350000 ;
      RECT 1016.500000 335.650000 1058.500000 336.350000 ;
      RECT 966.500000 335.650000 1008.500000 336.350000 ;
      RECT 916.500000 335.650000 958.500000 336.350000 ;
      RECT 866.500000 335.650000 908.500000 336.350000 ;
      RECT 816.500000 335.650000 858.500000 336.350000 ;
      RECT 766.500000 335.650000 808.500000 336.350000 ;
      RECT 716.500000 335.650000 758.500000 336.350000 ;
      RECT 666.500000 335.650000 708.500000 336.350000 ;
      RECT 616.500000 335.650000 658.500000 336.350000 ;
      RECT 566.500000 335.650000 608.500000 336.350000 ;
      RECT 516.500000 335.650000 558.500000 336.350000 ;
      RECT 466.500000 335.650000 508.500000 336.350000 ;
      RECT 416.500000 335.650000 458.500000 336.350000 ;
      RECT 366.500000 335.650000 408.500000 336.350000 ;
      RECT 316.500000 335.650000 358.500000 336.350000 ;
      RECT 266.500000 335.650000 308.500000 336.350000 ;
      RECT 216.500000 335.650000 258.500000 336.350000 ;
      RECT 166.500000 335.650000 208.500000 336.350000 ;
      RECT 116.500000 335.650000 158.500000 336.350000 ;
      RECT 66.500000 335.650000 108.500000 336.350000 ;
      RECT 29.500000 335.650000 58.500000 336.350000 ;
      RECT 0.000000 335.650000 16.500000 336.350000 ;
      RECT 1169.500000 334.350000 1170.500000 335.650000 ;
      RECT 1116.500000 334.350000 1149.500000 335.650000 ;
      RECT 1107.500000 334.350000 1108.500000 335.650000 ;
      RECT 1066.500000 334.350000 1099.500000 335.650000 ;
      RECT 1057.500000 334.350000 1058.500000 335.650000 ;
      RECT 1016.500000 334.350000 1049.500000 335.650000 ;
      RECT 1007.500000 334.350000 1008.500000 335.650000 ;
      RECT 966.500000 334.350000 999.500000 335.650000 ;
      RECT 957.500000 334.350000 958.500000 335.650000 ;
      RECT 916.500000 334.350000 949.500000 335.650000 ;
      RECT 907.500000 334.350000 908.500000 335.650000 ;
      RECT 866.500000 334.350000 899.500000 335.650000 ;
      RECT 857.500000 334.350000 858.500000 335.650000 ;
      RECT 816.500000 334.350000 849.500000 335.650000 ;
      RECT 807.500000 334.350000 808.500000 335.650000 ;
      RECT 766.500000 334.350000 799.500000 335.650000 ;
      RECT 757.500000 334.350000 758.500000 335.650000 ;
      RECT 716.500000 334.350000 749.500000 335.650000 ;
      RECT 707.500000 334.350000 708.500000 335.650000 ;
      RECT 666.500000 334.350000 699.500000 335.650000 ;
      RECT 657.500000 334.350000 658.500000 335.650000 ;
      RECT 616.500000 334.350000 649.500000 335.650000 ;
      RECT 607.500000 334.350000 608.500000 335.650000 ;
      RECT 566.500000 334.350000 599.500000 335.650000 ;
      RECT 557.500000 334.350000 558.500000 335.650000 ;
      RECT 516.500000 334.350000 549.500000 335.650000 ;
      RECT 507.500000 334.350000 508.500000 335.650000 ;
      RECT 466.500000 334.350000 499.500000 335.650000 ;
      RECT 457.500000 334.350000 458.500000 335.650000 ;
      RECT 416.500000 334.350000 449.500000 335.650000 ;
      RECT 407.500000 334.350000 408.500000 335.650000 ;
      RECT 366.500000 334.350000 399.500000 335.650000 ;
      RECT 357.500000 334.350000 358.500000 335.650000 ;
      RECT 316.500000 334.350000 349.500000 335.650000 ;
      RECT 307.500000 334.350000 308.500000 335.650000 ;
      RECT 266.500000 334.350000 299.500000 335.650000 ;
      RECT 257.500000 334.350000 258.500000 335.650000 ;
      RECT 216.500000 334.350000 249.500000 335.650000 ;
      RECT 207.500000 334.350000 208.500000 335.650000 ;
      RECT 166.500000 334.350000 199.500000 335.650000 ;
      RECT 157.500000 334.350000 158.500000 335.650000 ;
      RECT 116.500000 334.350000 149.500000 335.650000 ;
      RECT 107.500000 334.350000 108.500000 335.650000 ;
      RECT 66.500000 334.350000 99.500000 335.650000 ;
      RECT 57.500000 334.350000 58.500000 335.650000 ;
      RECT 29.500000 334.350000 49.500000 335.650000 ;
      RECT 15.500000 334.350000 16.500000 335.650000 ;
      RECT 1157.500000 333.650000 1170.500000 334.350000 ;
      RECT 1107.500000 333.650000 1149.500000 334.350000 ;
      RECT 1057.500000 333.650000 1099.500000 334.350000 ;
      RECT 1007.500000 333.650000 1049.500000 334.350000 ;
      RECT 957.500000 333.650000 999.500000 334.350000 ;
      RECT 907.500000 333.650000 949.500000 334.350000 ;
      RECT 857.500000 333.650000 899.500000 334.350000 ;
      RECT 807.500000 333.650000 849.500000 334.350000 ;
      RECT 757.500000 333.650000 799.500000 334.350000 ;
      RECT 707.500000 333.650000 749.500000 334.350000 ;
      RECT 657.500000 333.650000 699.500000 334.350000 ;
      RECT 607.500000 333.650000 649.500000 334.350000 ;
      RECT 557.500000 333.650000 599.500000 334.350000 ;
      RECT 507.500000 333.650000 549.500000 334.350000 ;
      RECT 457.500000 333.650000 499.500000 334.350000 ;
      RECT 407.500000 333.650000 449.500000 334.350000 ;
      RECT 357.500000 333.650000 399.500000 334.350000 ;
      RECT 307.500000 333.650000 349.500000 334.350000 ;
      RECT 257.500000 333.650000 299.500000 334.350000 ;
      RECT 207.500000 333.650000 249.500000 334.350000 ;
      RECT 157.500000 333.650000 199.500000 334.350000 ;
      RECT 107.500000 333.650000 149.500000 334.350000 ;
      RECT 57.500000 333.650000 99.500000 334.350000 ;
      RECT 15.500000 333.650000 49.500000 334.350000 ;
      RECT 1183.500000 332.350000 1186.000000 335.650000 ;
      RECT 1169.500000 332.350000 1170.500000 333.650000 ;
      RECT 1116.500000 332.350000 1149.500000 333.650000 ;
      RECT 1107.500000 332.350000 1108.500000 333.650000 ;
      RECT 1066.500000 332.350000 1099.500000 333.650000 ;
      RECT 1057.500000 332.350000 1058.500000 333.650000 ;
      RECT 1016.500000 332.350000 1049.500000 333.650000 ;
      RECT 1007.500000 332.350000 1008.500000 333.650000 ;
      RECT 966.500000 332.350000 999.500000 333.650000 ;
      RECT 957.500000 332.350000 958.500000 333.650000 ;
      RECT 916.500000 332.350000 949.500000 333.650000 ;
      RECT 907.500000 332.350000 908.500000 333.650000 ;
      RECT 866.500000 332.350000 899.500000 333.650000 ;
      RECT 857.500000 332.350000 858.500000 333.650000 ;
      RECT 816.500000 332.350000 849.500000 333.650000 ;
      RECT 807.500000 332.350000 808.500000 333.650000 ;
      RECT 766.500000 332.350000 799.500000 333.650000 ;
      RECT 757.500000 332.350000 758.500000 333.650000 ;
      RECT 716.500000 332.350000 749.500000 333.650000 ;
      RECT 707.500000 332.350000 708.500000 333.650000 ;
      RECT 666.500000 332.350000 699.500000 333.650000 ;
      RECT 657.500000 332.350000 658.500000 333.650000 ;
      RECT 616.500000 332.350000 649.500000 333.650000 ;
      RECT 607.500000 332.350000 608.500000 333.650000 ;
      RECT 566.500000 332.350000 599.500000 333.650000 ;
      RECT 557.500000 332.350000 558.500000 333.650000 ;
      RECT 516.500000 332.350000 549.500000 333.650000 ;
      RECT 507.500000 332.350000 508.500000 333.650000 ;
      RECT 466.500000 332.350000 499.500000 333.650000 ;
      RECT 457.500000 332.350000 458.500000 333.650000 ;
      RECT 416.500000 332.350000 449.500000 333.650000 ;
      RECT 407.500000 332.350000 408.500000 333.650000 ;
      RECT 366.500000 332.350000 399.500000 333.650000 ;
      RECT 357.500000 332.350000 358.500000 333.650000 ;
      RECT 316.500000 332.350000 349.500000 333.650000 ;
      RECT 307.500000 332.350000 308.500000 333.650000 ;
      RECT 266.500000 332.350000 299.500000 333.650000 ;
      RECT 257.500000 332.350000 258.500000 333.650000 ;
      RECT 216.500000 332.350000 249.500000 333.650000 ;
      RECT 207.500000 332.350000 208.500000 333.650000 ;
      RECT 166.500000 332.350000 199.500000 333.650000 ;
      RECT 157.500000 332.350000 158.500000 333.650000 ;
      RECT 116.500000 332.350000 149.500000 333.650000 ;
      RECT 107.500000 332.350000 108.500000 333.650000 ;
      RECT 66.500000 332.350000 99.500000 333.650000 ;
      RECT 57.500000 332.350000 58.500000 333.650000 ;
      RECT 29.500000 332.350000 49.500000 333.650000 ;
      RECT 15.500000 332.350000 16.500000 333.650000 ;
      RECT 0.000000 332.350000 2.500000 335.650000 ;
      RECT 1169.500000 331.650000 1186.000000 332.350000 ;
      RECT 1116.500000 331.650000 1156.500000 332.350000 ;
      RECT 1066.500000 331.650000 1108.500000 332.350000 ;
      RECT 1016.500000 331.650000 1058.500000 332.350000 ;
      RECT 966.500000 331.650000 1008.500000 332.350000 ;
      RECT 916.500000 331.650000 958.500000 332.350000 ;
      RECT 866.500000 331.650000 908.500000 332.350000 ;
      RECT 816.500000 331.650000 858.500000 332.350000 ;
      RECT 766.500000 331.650000 808.500000 332.350000 ;
      RECT 716.500000 331.650000 758.500000 332.350000 ;
      RECT 666.500000 331.650000 708.500000 332.350000 ;
      RECT 616.500000 331.650000 658.500000 332.350000 ;
      RECT 566.500000 331.650000 608.500000 332.350000 ;
      RECT 516.500000 331.650000 558.500000 332.350000 ;
      RECT 466.500000 331.650000 508.500000 332.350000 ;
      RECT 416.500000 331.650000 458.500000 332.350000 ;
      RECT 366.500000 331.650000 408.500000 332.350000 ;
      RECT 316.500000 331.650000 358.500000 332.350000 ;
      RECT 266.500000 331.650000 308.500000 332.350000 ;
      RECT 216.500000 331.650000 258.500000 332.350000 ;
      RECT 166.500000 331.650000 208.500000 332.350000 ;
      RECT 116.500000 331.650000 158.500000 332.350000 ;
      RECT 66.500000 331.650000 108.500000 332.350000 ;
      RECT 29.500000 331.650000 58.500000 332.350000 ;
      RECT 0.000000 331.650000 16.500000 332.350000 ;
      RECT 1169.500000 330.350000 1170.500000 331.650000 ;
      RECT 1116.500000 330.350000 1149.500000 331.650000 ;
      RECT 1107.500000 330.350000 1108.500000 331.650000 ;
      RECT 1066.500000 330.350000 1099.500000 331.650000 ;
      RECT 1057.500000 330.350000 1058.500000 331.650000 ;
      RECT 1016.500000 330.350000 1049.500000 331.650000 ;
      RECT 1007.500000 330.350000 1008.500000 331.650000 ;
      RECT 966.500000 330.350000 999.500000 331.650000 ;
      RECT 957.500000 330.350000 958.500000 331.650000 ;
      RECT 916.500000 330.350000 949.500000 331.650000 ;
      RECT 907.500000 330.350000 908.500000 331.650000 ;
      RECT 866.500000 330.350000 899.500000 331.650000 ;
      RECT 857.500000 330.350000 858.500000 331.650000 ;
      RECT 816.500000 330.350000 849.500000 331.650000 ;
      RECT 807.500000 330.350000 808.500000 331.650000 ;
      RECT 766.500000 330.350000 799.500000 331.650000 ;
      RECT 757.500000 330.350000 758.500000 331.650000 ;
      RECT 716.500000 330.350000 749.500000 331.650000 ;
      RECT 707.500000 330.350000 708.500000 331.650000 ;
      RECT 666.500000 330.350000 699.500000 331.650000 ;
      RECT 657.500000 330.350000 658.500000 331.650000 ;
      RECT 616.500000 330.350000 649.500000 331.650000 ;
      RECT 607.500000 330.350000 608.500000 331.650000 ;
      RECT 566.500000 330.350000 599.500000 331.650000 ;
      RECT 557.500000 330.350000 558.500000 331.650000 ;
      RECT 516.500000 330.350000 549.500000 331.650000 ;
      RECT 507.500000 330.350000 508.500000 331.650000 ;
      RECT 466.500000 330.350000 499.500000 331.650000 ;
      RECT 457.500000 330.350000 458.500000 331.650000 ;
      RECT 416.500000 330.350000 449.500000 331.650000 ;
      RECT 407.500000 330.350000 408.500000 331.650000 ;
      RECT 366.500000 330.350000 399.500000 331.650000 ;
      RECT 357.500000 330.350000 358.500000 331.650000 ;
      RECT 316.500000 330.350000 349.500000 331.650000 ;
      RECT 307.500000 330.350000 308.500000 331.650000 ;
      RECT 266.500000 330.350000 299.500000 331.650000 ;
      RECT 257.500000 330.350000 258.500000 331.650000 ;
      RECT 216.500000 330.350000 249.500000 331.650000 ;
      RECT 207.500000 330.350000 208.500000 331.650000 ;
      RECT 166.500000 330.350000 199.500000 331.650000 ;
      RECT 157.500000 330.350000 158.500000 331.650000 ;
      RECT 116.500000 330.350000 149.500000 331.650000 ;
      RECT 107.500000 330.350000 108.500000 331.650000 ;
      RECT 66.500000 330.350000 99.500000 331.650000 ;
      RECT 57.500000 330.350000 58.500000 331.650000 ;
      RECT 29.500000 330.350000 49.500000 331.650000 ;
      RECT 15.500000 330.350000 16.500000 331.650000 ;
      RECT 1157.500000 329.650000 1170.500000 330.350000 ;
      RECT 1107.500000 329.650000 1149.500000 330.350000 ;
      RECT 1057.500000 329.650000 1099.500000 330.350000 ;
      RECT 1007.500000 329.650000 1049.500000 330.350000 ;
      RECT 957.500000 329.650000 999.500000 330.350000 ;
      RECT 907.500000 329.650000 949.500000 330.350000 ;
      RECT 857.500000 329.650000 899.500000 330.350000 ;
      RECT 807.500000 329.650000 849.500000 330.350000 ;
      RECT 757.500000 329.650000 799.500000 330.350000 ;
      RECT 707.500000 329.650000 749.500000 330.350000 ;
      RECT 657.500000 329.650000 699.500000 330.350000 ;
      RECT 607.500000 329.650000 649.500000 330.350000 ;
      RECT 557.500000 329.650000 599.500000 330.350000 ;
      RECT 507.500000 329.650000 549.500000 330.350000 ;
      RECT 457.500000 329.650000 499.500000 330.350000 ;
      RECT 407.500000 329.650000 449.500000 330.350000 ;
      RECT 357.500000 329.650000 399.500000 330.350000 ;
      RECT 307.500000 329.650000 349.500000 330.350000 ;
      RECT 257.500000 329.650000 299.500000 330.350000 ;
      RECT 207.500000 329.650000 249.500000 330.350000 ;
      RECT 157.500000 329.650000 199.500000 330.350000 ;
      RECT 107.500000 329.650000 149.500000 330.350000 ;
      RECT 57.500000 329.650000 99.500000 330.350000 ;
      RECT 15.500000 329.650000 49.500000 330.350000 ;
      RECT 1183.500000 328.350000 1186.000000 331.650000 ;
      RECT 1169.500000 328.350000 1170.500000 329.650000 ;
      RECT 1116.500000 328.350000 1149.500000 329.650000 ;
      RECT 1107.500000 328.350000 1108.500000 329.650000 ;
      RECT 1066.500000 328.350000 1099.500000 329.650000 ;
      RECT 1057.500000 328.350000 1058.500000 329.650000 ;
      RECT 1016.500000 328.350000 1049.500000 329.650000 ;
      RECT 1007.500000 328.350000 1008.500000 329.650000 ;
      RECT 966.500000 328.350000 999.500000 329.650000 ;
      RECT 957.500000 328.350000 958.500000 329.650000 ;
      RECT 916.500000 328.350000 949.500000 329.650000 ;
      RECT 907.500000 328.350000 908.500000 329.650000 ;
      RECT 866.500000 328.350000 899.500000 329.650000 ;
      RECT 857.500000 328.350000 858.500000 329.650000 ;
      RECT 816.500000 328.350000 849.500000 329.650000 ;
      RECT 807.500000 328.350000 808.500000 329.650000 ;
      RECT 766.500000 328.350000 799.500000 329.650000 ;
      RECT 757.500000 328.350000 758.500000 329.650000 ;
      RECT 716.500000 328.350000 749.500000 329.650000 ;
      RECT 707.500000 328.350000 708.500000 329.650000 ;
      RECT 666.500000 328.350000 699.500000 329.650000 ;
      RECT 657.500000 328.350000 658.500000 329.650000 ;
      RECT 616.500000 328.350000 649.500000 329.650000 ;
      RECT 607.500000 328.350000 608.500000 329.650000 ;
      RECT 566.500000 328.350000 599.500000 329.650000 ;
      RECT 557.500000 328.350000 558.500000 329.650000 ;
      RECT 516.500000 328.350000 549.500000 329.650000 ;
      RECT 507.500000 328.350000 508.500000 329.650000 ;
      RECT 466.500000 328.350000 499.500000 329.650000 ;
      RECT 457.500000 328.350000 458.500000 329.650000 ;
      RECT 416.500000 328.350000 449.500000 329.650000 ;
      RECT 407.500000 328.350000 408.500000 329.650000 ;
      RECT 366.500000 328.350000 399.500000 329.650000 ;
      RECT 357.500000 328.350000 358.500000 329.650000 ;
      RECT 316.500000 328.350000 349.500000 329.650000 ;
      RECT 307.500000 328.350000 308.500000 329.650000 ;
      RECT 266.500000 328.350000 299.500000 329.650000 ;
      RECT 257.500000 328.350000 258.500000 329.650000 ;
      RECT 216.500000 328.350000 249.500000 329.650000 ;
      RECT 207.500000 328.350000 208.500000 329.650000 ;
      RECT 166.500000 328.350000 199.500000 329.650000 ;
      RECT 157.500000 328.350000 158.500000 329.650000 ;
      RECT 116.500000 328.350000 149.500000 329.650000 ;
      RECT 107.500000 328.350000 108.500000 329.650000 ;
      RECT 66.500000 328.350000 99.500000 329.650000 ;
      RECT 57.500000 328.350000 58.500000 329.650000 ;
      RECT 29.500000 328.350000 49.500000 329.650000 ;
      RECT 15.500000 328.350000 16.500000 329.650000 ;
      RECT 0.000000 328.350000 2.500000 331.650000 ;
      RECT 1169.500000 327.650000 1186.000000 328.350000 ;
      RECT 1116.500000 327.650000 1156.500000 328.350000 ;
      RECT 1066.500000 327.650000 1108.500000 328.350000 ;
      RECT 1016.500000 327.650000 1058.500000 328.350000 ;
      RECT 966.500000 327.650000 1008.500000 328.350000 ;
      RECT 916.500000 327.650000 958.500000 328.350000 ;
      RECT 866.500000 327.650000 908.500000 328.350000 ;
      RECT 816.500000 327.650000 858.500000 328.350000 ;
      RECT 766.500000 327.650000 808.500000 328.350000 ;
      RECT 716.500000 327.650000 758.500000 328.350000 ;
      RECT 666.500000 327.650000 708.500000 328.350000 ;
      RECT 616.500000 327.650000 658.500000 328.350000 ;
      RECT 566.500000 327.650000 608.500000 328.350000 ;
      RECT 516.500000 327.650000 558.500000 328.350000 ;
      RECT 466.500000 327.650000 508.500000 328.350000 ;
      RECT 416.500000 327.650000 458.500000 328.350000 ;
      RECT 366.500000 327.650000 408.500000 328.350000 ;
      RECT 316.500000 327.650000 358.500000 328.350000 ;
      RECT 266.500000 327.650000 308.500000 328.350000 ;
      RECT 216.500000 327.650000 258.500000 328.350000 ;
      RECT 166.500000 327.650000 208.500000 328.350000 ;
      RECT 116.500000 327.650000 158.500000 328.350000 ;
      RECT 66.500000 327.650000 108.500000 328.350000 ;
      RECT 29.500000 327.650000 58.500000 328.350000 ;
      RECT 0.000000 327.650000 16.500000 328.350000 ;
      RECT 1169.500000 326.350000 1170.500000 327.650000 ;
      RECT 1116.500000 326.350000 1149.500000 327.650000 ;
      RECT 1107.500000 326.350000 1108.500000 327.650000 ;
      RECT 1066.500000 326.350000 1099.500000 327.650000 ;
      RECT 1057.500000 326.350000 1058.500000 327.650000 ;
      RECT 1016.500000 326.350000 1049.500000 327.650000 ;
      RECT 1007.500000 326.350000 1008.500000 327.650000 ;
      RECT 966.500000 326.350000 999.500000 327.650000 ;
      RECT 957.500000 326.350000 958.500000 327.650000 ;
      RECT 916.500000 326.350000 949.500000 327.650000 ;
      RECT 907.500000 326.350000 908.500000 327.650000 ;
      RECT 866.500000 326.350000 899.500000 327.650000 ;
      RECT 857.500000 326.350000 858.500000 327.650000 ;
      RECT 816.500000 326.350000 849.500000 327.650000 ;
      RECT 807.500000 326.350000 808.500000 327.650000 ;
      RECT 766.500000 326.350000 799.500000 327.650000 ;
      RECT 757.500000 326.350000 758.500000 327.650000 ;
      RECT 716.500000 326.350000 749.500000 327.650000 ;
      RECT 707.500000 326.350000 708.500000 327.650000 ;
      RECT 666.500000 326.350000 699.500000 327.650000 ;
      RECT 657.500000 326.350000 658.500000 327.650000 ;
      RECT 616.500000 326.350000 649.500000 327.650000 ;
      RECT 607.500000 326.350000 608.500000 327.650000 ;
      RECT 566.500000 326.350000 599.500000 327.650000 ;
      RECT 557.500000 326.350000 558.500000 327.650000 ;
      RECT 516.500000 326.350000 549.500000 327.650000 ;
      RECT 507.500000 326.350000 508.500000 327.650000 ;
      RECT 466.500000 326.350000 499.500000 327.650000 ;
      RECT 457.500000 326.350000 458.500000 327.650000 ;
      RECT 416.500000 326.350000 449.500000 327.650000 ;
      RECT 407.500000 326.350000 408.500000 327.650000 ;
      RECT 366.500000 326.350000 399.500000 327.650000 ;
      RECT 357.500000 326.350000 358.500000 327.650000 ;
      RECT 316.500000 326.350000 349.500000 327.650000 ;
      RECT 307.500000 326.350000 308.500000 327.650000 ;
      RECT 266.500000 326.350000 299.500000 327.650000 ;
      RECT 257.500000 326.350000 258.500000 327.650000 ;
      RECT 216.500000 326.350000 249.500000 327.650000 ;
      RECT 207.500000 326.350000 208.500000 327.650000 ;
      RECT 166.500000 326.350000 199.500000 327.650000 ;
      RECT 157.500000 326.350000 158.500000 327.650000 ;
      RECT 116.500000 326.350000 149.500000 327.650000 ;
      RECT 107.500000 326.350000 108.500000 327.650000 ;
      RECT 66.500000 326.350000 99.500000 327.650000 ;
      RECT 57.500000 326.350000 58.500000 327.650000 ;
      RECT 29.500000 326.350000 49.500000 327.650000 ;
      RECT 15.500000 326.350000 16.500000 327.650000 ;
      RECT 1157.500000 325.650000 1170.500000 326.350000 ;
      RECT 1107.500000 325.650000 1149.500000 326.350000 ;
      RECT 1057.500000 325.650000 1099.500000 326.350000 ;
      RECT 1007.500000 325.650000 1049.500000 326.350000 ;
      RECT 957.500000 325.650000 999.500000 326.350000 ;
      RECT 907.500000 325.650000 949.500000 326.350000 ;
      RECT 857.500000 325.650000 899.500000 326.350000 ;
      RECT 807.500000 325.650000 849.500000 326.350000 ;
      RECT 757.500000 325.650000 799.500000 326.350000 ;
      RECT 707.500000 325.650000 749.500000 326.350000 ;
      RECT 657.500000 325.650000 699.500000 326.350000 ;
      RECT 607.500000 325.650000 649.500000 326.350000 ;
      RECT 557.500000 325.650000 599.500000 326.350000 ;
      RECT 507.500000 325.650000 549.500000 326.350000 ;
      RECT 457.500000 325.650000 499.500000 326.350000 ;
      RECT 407.500000 325.650000 449.500000 326.350000 ;
      RECT 357.500000 325.650000 399.500000 326.350000 ;
      RECT 307.500000 325.650000 349.500000 326.350000 ;
      RECT 257.500000 325.650000 299.500000 326.350000 ;
      RECT 207.500000 325.650000 249.500000 326.350000 ;
      RECT 157.500000 325.650000 199.500000 326.350000 ;
      RECT 107.500000 325.650000 149.500000 326.350000 ;
      RECT 57.500000 325.650000 99.500000 326.350000 ;
      RECT 15.500000 325.650000 49.500000 326.350000 ;
      RECT 1183.500000 324.350000 1186.000000 327.650000 ;
      RECT 1169.500000 324.350000 1170.500000 325.650000 ;
      RECT 1116.500000 324.350000 1149.500000 325.650000 ;
      RECT 1107.500000 324.350000 1108.500000 325.650000 ;
      RECT 1066.500000 324.350000 1099.500000 325.650000 ;
      RECT 1057.500000 324.350000 1058.500000 325.650000 ;
      RECT 1016.500000 324.350000 1049.500000 325.650000 ;
      RECT 1007.500000 324.350000 1008.500000 325.650000 ;
      RECT 966.500000 324.350000 999.500000 325.650000 ;
      RECT 957.500000 324.350000 958.500000 325.650000 ;
      RECT 916.500000 324.350000 949.500000 325.650000 ;
      RECT 907.500000 324.350000 908.500000 325.650000 ;
      RECT 866.500000 324.350000 899.500000 325.650000 ;
      RECT 857.500000 324.350000 858.500000 325.650000 ;
      RECT 816.500000 324.350000 849.500000 325.650000 ;
      RECT 807.500000 324.350000 808.500000 325.650000 ;
      RECT 766.500000 324.350000 799.500000 325.650000 ;
      RECT 757.500000 324.350000 758.500000 325.650000 ;
      RECT 716.500000 324.350000 749.500000 325.650000 ;
      RECT 707.500000 324.350000 708.500000 325.650000 ;
      RECT 666.500000 324.350000 699.500000 325.650000 ;
      RECT 657.500000 324.350000 658.500000 325.650000 ;
      RECT 616.500000 324.350000 649.500000 325.650000 ;
      RECT 607.500000 324.350000 608.500000 325.650000 ;
      RECT 566.500000 324.350000 599.500000 325.650000 ;
      RECT 557.500000 324.350000 558.500000 325.650000 ;
      RECT 516.500000 324.350000 549.500000 325.650000 ;
      RECT 507.500000 324.350000 508.500000 325.650000 ;
      RECT 466.500000 324.350000 499.500000 325.650000 ;
      RECT 457.500000 324.350000 458.500000 325.650000 ;
      RECT 416.500000 324.350000 449.500000 325.650000 ;
      RECT 407.500000 324.350000 408.500000 325.650000 ;
      RECT 366.500000 324.350000 399.500000 325.650000 ;
      RECT 357.500000 324.350000 358.500000 325.650000 ;
      RECT 316.500000 324.350000 349.500000 325.650000 ;
      RECT 307.500000 324.350000 308.500000 325.650000 ;
      RECT 266.500000 324.350000 299.500000 325.650000 ;
      RECT 257.500000 324.350000 258.500000 325.650000 ;
      RECT 216.500000 324.350000 249.500000 325.650000 ;
      RECT 207.500000 324.350000 208.500000 325.650000 ;
      RECT 166.500000 324.350000 199.500000 325.650000 ;
      RECT 157.500000 324.350000 158.500000 325.650000 ;
      RECT 116.500000 324.350000 149.500000 325.650000 ;
      RECT 107.500000 324.350000 108.500000 325.650000 ;
      RECT 66.500000 324.350000 99.500000 325.650000 ;
      RECT 57.500000 324.350000 58.500000 325.650000 ;
      RECT 29.500000 324.350000 49.500000 325.650000 ;
      RECT 15.500000 324.350000 16.500000 325.650000 ;
      RECT 0.000000 324.350000 2.500000 327.650000 ;
      RECT 1169.500000 323.650000 1186.000000 324.350000 ;
      RECT 1116.500000 323.650000 1156.500000 324.350000 ;
      RECT 1066.500000 323.650000 1108.500000 324.350000 ;
      RECT 1016.500000 323.650000 1058.500000 324.350000 ;
      RECT 966.500000 323.650000 1008.500000 324.350000 ;
      RECT 916.500000 323.650000 958.500000 324.350000 ;
      RECT 866.500000 323.650000 908.500000 324.350000 ;
      RECT 816.500000 323.650000 858.500000 324.350000 ;
      RECT 766.500000 323.650000 808.500000 324.350000 ;
      RECT 716.500000 323.650000 758.500000 324.350000 ;
      RECT 666.500000 323.650000 708.500000 324.350000 ;
      RECT 616.500000 323.650000 658.500000 324.350000 ;
      RECT 566.500000 323.650000 608.500000 324.350000 ;
      RECT 516.500000 323.650000 558.500000 324.350000 ;
      RECT 466.500000 323.650000 508.500000 324.350000 ;
      RECT 416.500000 323.650000 458.500000 324.350000 ;
      RECT 366.500000 323.650000 408.500000 324.350000 ;
      RECT 316.500000 323.650000 358.500000 324.350000 ;
      RECT 266.500000 323.650000 308.500000 324.350000 ;
      RECT 216.500000 323.650000 258.500000 324.350000 ;
      RECT 166.500000 323.650000 208.500000 324.350000 ;
      RECT 116.500000 323.650000 158.500000 324.350000 ;
      RECT 66.500000 323.650000 108.500000 324.350000 ;
      RECT 29.500000 323.650000 58.500000 324.350000 ;
      RECT 0.000000 323.650000 16.500000 324.350000 ;
      RECT 1169.500000 322.350000 1170.500000 323.650000 ;
      RECT 1116.500000 322.350000 1149.500000 323.650000 ;
      RECT 1107.500000 322.350000 1108.500000 323.650000 ;
      RECT 1066.500000 322.350000 1099.500000 323.650000 ;
      RECT 1057.500000 322.350000 1058.500000 323.650000 ;
      RECT 1016.500000 322.350000 1049.500000 323.650000 ;
      RECT 1007.500000 322.350000 1008.500000 323.650000 ;
      RECT 966.500000 322.350000 999.500000 323.650000 ;
      RECT 957.500000 322.350000 958.500000 323.650000 ;
      RECT 916.500000 322.350000 949.500000 323.650000 ;
      RECT 907.500000 322.350000 908.500000 323.650000 ;
      RECT 866.500000 322.350000 899.500000 323.650000 ;
      RECT 857.500000 322.350000 858.500000 323.650000 ;
      RECT 816.500000 322.350000 849.500000 323.650000 ;
      RECT 807.500000 322.350000 808.500000 323.650000 ;
      RECT 766.500000 322.350000 799.500000 323.650000 ;
      RECT 757.500000 322.350000 758.500000 323.650000 ;
      RECT 716.500000 322.350000 749.500000 323.650000 ;
      RECT 707.500000 322.350000 708.500000 323.650000 ;
      RECT 666.500000 322.350000 699.500000 323.650000 ;
      RECT 657.500000 322.350000 658.500000 323.650000 ;
      RECT 616.500000 322.350000 649.500000 323.650000 ;
      RECT 607.500000 322.350000 608.500000 323.650000 ;
      RECT 566.500000 322.350000 599.500000 323.650000 ;
      RECT 557.500000 322.350000 558.500000 323.650000 ;
      RECT 516.500000 322.350000 549.500000 323.650000 ;
      RECT 507.500000 322.350000 508.500000 323.650000 ;
      RECT 466.500000 322.350000 499.500000 323.650000 ;
      RECT 457.500000 322.350000 458.500000 323.650000 ;
      RECT 416.500000 322.350000 449.500000 323.650000 ;
      RECT 407.500000 322.350000 408.500000 323.650000 ;
      RECT 366.500000 322.350000 399.500000 323.650000 ;
      RECT 357.500000 322.350000 358.500000 323.650000 ;
      RECT 316.500000 322.350000 349.500000 323.650000 ;
      RECT 307.500000 322.350000 308.500000 323.650000 ;
      RECT 266.500000 322.350000 299.500000 323.650000 ;
      RECT 257.500000 322.350000 258.500000 323.650000 ;
      RECT 216.500000 322.350000 249.500000 323.650000 ;
      RECT 207.500000 322.350000 208.500000 323.650000 ;
      RECT 166.500000 322.350000 199.500000 323.650000 ;
      RECT 157.500000 322.350000 158.500000 323.650000 ;
      RECT 116.500000 322.350000 149.500000 323.650000 ;
      RECT 107.500000 322.350000 108.500000 323.650000 ;
      RECT 66.500000 322.350000 99.500000 323.650000 ;
      RECT 57.500000 322.350000 58.500000 323.650000 ;
      RECT 29.500000 322.350000 49.500000 323.650000 ;
      RECT 15.500000 322.350000 16.500000 323.650000 ;
      RECT 1157.500000 321.650000 1170.500000 322.350000 ;
      RECT 1107.500000 321.650000 1149.500000 322.350000 ;
      RECT 1057.500000 321.650000 1099.500000 322.350000 ;
      RECT 1007.500000 321.650000 1049.500000 322.350000 ;
      RECT 957.500000 321.650000 999.500000 322.350000 ;
      RECT 907.500000 321.650000 949.500000 322.350000 ;
      RECT 857.500000 321.650000 899.500000 322.350000 ;
      RECT 807.500000 321.650000 849.500000 322.350000 ;
      RECT 757.500000 321.650000 799.500000 322.350000 ;
      RECT 707.500000 321.650000 749.500000 322.350000 ;
      RECT 657.500000 321.650000 699.500000 322.350000 ;
      RECT 607.500000 321.650000 649.500000 322.350000 ;
      RECT 557.500000 321.650000 599.500000 322.350000 ;
      RECT 507.500000 321.650000 549.500000 322.350000 ;
      RECT 457.500000 321.650000 499.500000 322.350000 ;
      RECT 407.500000 321.650000 449.500000 322.350000 ;
      RECT 357.500000 321.650000 399.500000 322.350000 ;
      RECT 307.500000 321.650000 349.500000 322.350000 ;
      RECT 257.500000 321.650000 299.500000 322.350000 ;
      RECT 207.500000 321.650000 249.500000 322.350000 ;
      RECT 157.500000 321.650000 199.500000 322.350000 ;
      RECT 107.500000 321.650000 149.500000 322.350000 ;
      RECT 57.500000 321.650000 99.500000 322.350000 ;
      RECT 15.500000 321.650000 49.500000 322.350000 ;
      RECT 1183.500000 320.350000 1186.000000 323.650000 ;
      RECT 1169.500000 320.350000 1170.500000 321.650000 ;
      RECT 1116.500000 320.350000 1149.500000 321.650000 ;
      RECT 1107.500000 320.350000 1108.500000 321.650000 ;
      RECT 1066.500000 320.350000 1099.500000 321.650000 ;
      RECT 1057.500000 320.350000 1058.500000 321.650000 ;
      RECT 1016.500000 320.350000 1049.500000 321.650000 ;
      RECT 1007.500000 320.350000 1008.500000 321.650000 ;
      RECT 966.500000 320.350000 999.500000 321.650000 ;
      RECT 957.500000 320.350000 958.500000 321.650000 ;
      RECT 916.500000 320.350000 949.500000 321.650000 ;
      RECT 907.500000 320.350000 908.500000 321.650000 ;
      RECT 866.500000 320.350000 899.500000 321.650000 ;
      RECT 857.500000 320.350000 858.500000 321.650000 ;
      RECT 816.500000 320.350000 849.500000 321.650000 ;
      RECT 807.500000 320.350000 808.500000 321.650000 ;
      RECT 766.500000 320.350000 799.500000 321.650000 ;
      RECT 757.500000 320.350000 758.500000 321.650000 ;
      RECT 716.500000 320.350000 749.500000 321.650000 ;
      RECT 707.500000 320.350000 708.500000 321.650000 ;
      RECT 666.500000 320.350000 699.500000 321.650000 ;
      RECT 657.500000 320.350000 658.500000 321.650000 ;
      RECT 616.500000 320.350000 649.500000 321.650000 ;
      RECT 607.500000 320.350000 608.500000 321.650000 ;
      RECT 566.500000 320.350000 599.500000 321.650000 ;
      RECT 557.500000 320.350000 558.500000 321.650000 ;
      RECT 516.500000 320.350000 549.500000 321.650000 ;
      RECT 507.500000 320.350000 508.500000 321.650000 ;
      RECT 466.500000 320.350000 499.500000 321.650000 ;
      RECT 457.500000 320.350000 458.500000 321.650000 ;
      RECT 416.500000 320.350000 449.500000 321.650000 ;
      RECT 407.500000 320.350000 408.500000 321.650000 ;
      RECT 366.500000 320.350000 399.500000 321.650000 ;
      RECT 357.500000 320.350000 358.500000 321.650000 ;
      RECT 316.500000 320.350000 349.500000 321.650000 ;
      RECT 307.500000 320.350000 308.500000 321.650000 ;
      RECT 266.500000 320.350000 299.500000 321.650000 ;
      RECT 257.500000 320.350000 258.500000 321.650000 ;
      RECT 216.500000 320.350000 249.500000 321.650000 ;
      RECT 207.500000 320.350000 208.500000 321.650000 ;
      RECT 166.500000 320.350000 199.500000 321.650000 ;
      RECT 157.500000 320.350000 158.500000 321.650000 ;
      RECT 116.500000 320.350000 149.500000 321.650000 ;
      RECT 107.500000 320.350000 108.500000 321.650000 ;
      RECT 66.500000 320.350000 99.500000 321.650000 ;
      RECT 57.500000 320.350000 58.500000 321.650000 ;
      RECT 29.500000 320.350000 49.500000 321.650000 ;
      RECT 15.500000 320.350000 16.500000 321.650000 ;
      RECT 0.000000 320.350000 2.500000 323.650000 ;
      RECT 1169.500000 319.650000 1186.000000 320.350000 ;
      RECT 1116.500000 319.650000 1156.500000 320.350000 ;
      RECT 1066.500000 319.650000 1108.500000 320.350000 ;
      RECT 1016.500000 319.650000 1058.500000 320.350000 ;
      RECT 966.500000 319.650000 1008.500000 320.350000 ;
      RECT 916.500000 319.650000 958.500000 320.350000 ;
      RECT 866.500000 319.650000 908.500000 320.350000 ;
      RECT 816.500000 319.650000 858.500000 320.350000 ;
      RECT 766.500000 319.650000 808.500000 320.350000 ;
      RECT 716.500000 319.650000 758.500000 320.350000 ;
      RECT 666.500000 319.650000 708.500000 320.350000 ;
      RECT 616.500000 319.650000 658.500000 320.350000 ;
      RECT 566.500000 319.650000 608.500000 320.350000 ;
      RECT 516.500000 319.650000 558.500000 320.350000 ;
      RECT 466.500000 319.650000 508.500000 320.350000 ;
      RECT 366.500000 319.650000 408.500000 320.350000 ;
      RECT 316.500000 319.650000 358.500000 320.350000 ;
      RECT 266.500000 319.650000 308.500000 320.350000 ;
      RECT 216.500000 319.650000 258.500000 320.350000 ;
      RECT 166.500000 319.650000 208.500000 320.350000 ;
      RECT 116.500000 319.650000 158.500000 320.350000 ;
      RECT 66.500000 319.650000 108.500000 320.350000 ;
      RECT 29.500000 319.650000 58.500000 320.350000 ;
      RECT 0.000000 319.650000 16.500000 320.350000 ;
      RECT 1169.500000 318.350000 1170.500000 319.650000 ;
      RECT 1116.500000 318.350000 1149.500000 319.650000 ;
      RECT 1107.500000 318.350000 1108.500000 319.650000 ;
      RECT 1066.500000 318.350000 1099.500000 319.650000 ;
      RECT 1057.500000 318.350000 1058.500000 319.650000 ;
      RECT 1016.500000 318.350000 1049.500000 319.650000 ;
      RECT 1007.500000 318.350000 1008.500000 319.650000 ;
      RECT 966.500000 318.350000 999.500000 319.650000 ;
      RECT 957.500000 318.350000 958.500000 319.650000 ;
      RECT 916.500000 318.350000 949.500000 319.650000 ;
      RECT 907.500000 318.350000 908.500000 319.650000 ;
      RECT 866.500000 318.350000 899.500000 319.650000 ;
      RECT 857.500000 318.350000 858.500000 319.650000 ;
      RECT 816.500000 318.350000 849.500000 319.650000 ;
      RECT 807.500000 318.350000 808.500000 319.650000 ;
      RECT 766.500000 318.350000 799.500000 319.650000 ;
      RECT 757.500000 318.350000 758.500000 319.650000 ;
      RECT 716.500000 318.350000 749.500000 319.650000 ;
      RECT 707.500000 318.350000 708.500000 319.650000 ;
      RECT 666.500000 318.350000 699.500000 319.650000 ;
      RECT 657.500000 318.350000 658.500000 319.650000 ;
      RECT 616.500000 318.350000 649.500000 319.650000 ;
      RECT 607.500000 318.350000 608.500000 319.650000 ;
      RECT 566.500000 318.350000 599.500000 319.650000 ;
      RECT 557.500000 318.350000 558.500000 319.650000 ;
      RECT 516.500000 318.350000 549.500000 319.650000 ;
      RECT 507.500000 318.350000 508.500000 319.650000 ;
      RECT 466.500000 318.350000 499.500000 319.650000 ;
      RECT 416.500000 318.350000 458.500000 320.350000 ;
      RECT 407.500000 318.350000 408.500000 319.650000 ;
      RECT 366.500000 318.350000 399.500000 319.650000 ;
      RECT 357.500000 318.350000 358.500000 319.650000 ;
      RECT 316.500000 318.350000 349.500000 319.650000 ;
      RECT 307.500000 318.350000 308.500000 319.650000 ;
      RECT 266.500000 318.350000 299.500000 319.650000 ;
      RECT 257.500000 318.350000 258.500000 319.650000 ;
      RECT 216.500000 318.350000 249.500000 319.650000 ;
      RECT 207.500000 318.350000 208.500000 319.650000 ;
      RECT 166.500000 318.350000 199.500000 319.650000 ;
      RECT 157.500000 318.350000 158.500000 319.650000 ;
      RECT 116.500000 318.350000 149.500000 319.650000 ;
      RECT 107.500000 318.350000 108.500000 319.650000 ;
      RECT 66.500000 318.350000 99.500000 319.650000 ;
      RECT 57.500000 318.350000 58.500000 319.650000 ;
      RECT 29.500000 318.350000 49.500000 319.650000 ;
      RECT 15.500000 318.350000 16.500000 319.650000 ;
      RECT 1157.500000 317.650000 1170.500000 318.350000 ;
      RECT 1107.500000 317.650000 1149.500000 318.350000 ;
      RECT 1057.500000 317.650000 1099.500000 318.350000 ;
      RECT 1007.500000 317.650000 1049.500000 318.350000 ;
      RECT 957.500000 317.650000 999.500000 318.350000 ;
      RECT 907.500000 317.650000 949.500000 318.350000 ;
      RECT 857.500000 317.650000 899.500000 318.350000 ;
      RECT 807.500000 317.650000 849.500000 318.350000 ;
      RECT 757.500000 317.650000 799.500000 318.350000 ;
      RECT 707.500000 317.650000 749.500000 318.350000 ;
      RECT 657.500000 317.650000 699.500000 318.350000 ;
      RECT 607.500000 317.650000 649.500000 318.350000 ;
      RECT 557.500000 317.650000 599.500000 318.350000 ;
      RECT 507.500000 317.650000 549.500000 318.350000 ;
      RECT 407.500000 317.650000 499.500000 318.350000 ;
      RECT 357.500000 317.650000 399.500000 318.350000 ;
      RECT 307.500000 317.650000 349.500000 318.350000 ;
      RECT 257.500000 317.650000 299.500000 318.350000 ;
      RECT 207.500000 317.650000 249.500000 318.350000 ;
      RECT 157.500000 317.650000 199.500000 318.350000 ;
      RECT 107.500000 317.650000 149.500000 318.350000 ;
      RECT 57.500000 317.650000 99.500000 318.350000 ;
      RECT 15.500000 317.650000 49.500000 318.350000 ;
      RECT 1183.500000 316.350000 1186.000000 319.650000 ;
      RECT 1169.500000 316.350000 1170.500000 317.650000 ;
      RECT 1116.500000 316.350000 1149.500000 317.650000 ;
      RECT 1107.500000 316.350000 1108.500000 317.650000 ;
      RECT 1066.500000 316.350000 1099.500000 317.650000 ;
      RECT 1057.500000 316.350000 1058.500000 317.650000 ;
      RECT 1016.500000 316.350000 1049.500000 317.650000 ;
      RECT 1007.500000 316.350000 1008.500000 317.650000 ;
      RECT 966.500000 316.350000 999.500000 317.650000 ;
      RECT 957.500000 316.350000 958.500000 317.650000 ;
      RECT 916.500000 316.350000 949.500000 317.650000 ;
      RECT 907.500000 316.350000 908.500000 317.650000 ;
      RECT 866.500000 316.350000 899.500000 317.650000 ;
      RECT 857.500000 316.350000 858.500000 317.650000 ;
      RECT 816.500000 316.350000 849.500000 317.650000 ;
      RECT 807.500000 316.350000 808.500000 317.650000 ;
      RECT 766.500000 316.350000 799.500000 317.650000 ;
      RECT 757.500000 316.350000 758.500000 317.650000 ;
      RECT 716.500000 316.350000 749.500000 317.650000 ;
      RECT 707.500000 316.350000 708.500000 317.650000 ;
      RECT 666.500000 316.350000 699.500000 317.650000 ;
      RECT 657.500000 316.350000 658.500000 317.650000 ;
      RECT 616.500000 316.350000 649.500000 317.650000 ;
      RECT 607.500000 316.350000 608.500000 317.650000 ;
      RECT 566.500000 316.350000 599.500000 317.650000 ;
      RECT 557.500000 316.350000 558.500000 317.650000 ;
      RECT 516.500000 316.350000 549.500000 317.650000 ;
      RECT 507.500000 316.350000 508.500000 317.650000 ;
      RECT 416.500000 316.350000 499.500000 317.650000 ;
      RECT 407.500000 316.350000 408.500000 317.650000 ;
      RECT 366.500000 316.350000 399.500000 317.650000 ;
      RECT 357.500000 316.350000 358.500000 317.650000 ;
      RECT 316.500000 316.350000 349.500000 317.650000 ;
      RECT 307.500000 316.350000 308.500000 317.650000 ;
      RECT 266.500000 316.350000 299.500000 317.650000 ;
      RECT 257.500000 316.350000 258.500000 317.650000 ;
      RECT 216.500000 316.350000 249.500000 317.650000 ;
      RECT 207.500000 316.350000 208.500000 317.650000 ;
      RECT 166.500000 316.350000 199.500000 317.650000 ;
      RECT 157.500000 316.350000 158.500000 317.650000 ;
      RECT 116.500000 316.350000 149.500000 317.650000 ;
      RECT 107.500000 316.350000 108.500000 317.650000 ;
      RECT 66.500000 316.350000 99.500000 317.650000 ;
      RECT 57.500000 316.350000 58.500000 317.650000 ;
      RECT 29.500000 316.350000 49.500000 317.650000 ;
      RECT 15.500000 316.350000 16.500000 317.650000 ;
      RECT 0.000000 316.350000 2.500000 319.650000 ;
      RECT 1169.500000 315.650000 1186.000000 316.350000 ;
      RECT 1116.500000 315.650000 1156.500000 316.350000 ;
      RECT 1066.500000 315.650000 1108.500000 316.350000 ;
      RECT 1016.500000 315.650000 1058.500000 316.350000 ;
      RECT 966.500000 315.650000 1008.500000 316.350000 ;
      RECT 916.500000 315.650000 958.500000 316.350000 ;
      RECT 866.500000 315.650000 908.500000 316.350000 ;
      RECT 816.500000 315.650000 858.500000 316.350000 ;
      RECT 766.500000 315.650000 808.500000 316.350000 ;
      RECT 716.500000 315.650000 758.500000 316.350000 ;
      RECT 666.500000 315.650000 708.500000 316.350000 ;
      RECT 616.500000 315.650000 658.500000 316.350000 ;
      RECT 566.500000 315.650000 608.500000 316.350000 ;
      RECT 516.500000 315.650000 558.500000 316.350000 ;
      RECT 416.500000 315.650000 508.500000 316.350000 ;
      RECT 366.500000 315.650000 408.500000 316.350000 ;
      RECT 316.500000 315.650000 358.500000 316.350000 ;
      RECT 266.500000 315.650000 308.500000 316.350000 ;
      RECT 216.500000 315.650000 258.500000 316.350000 ;
      RECT 166.500000 315.650000 208.500000 316.350000 ;
      RECT 116.500000 315.650000 158.500000 316.350000 ;
      RECT 66.500000 315.650000 108.500000 316.350000 ;
      RECT 29.500000 315.650000 58.500000 316.350000 ;
      RECT 0.000000 315.650000 16.500000 316.350000 ;
      RECT 1169.500000 314.350000 1170.500000 315.650000 ;
      RECT 1116.500000 314.350000 1149.500000 315.650000 ;
      RECT 1107.500000 314.350000 1108.500000 315.650000 ;
      RECT 1066.500000 314.350000 1099.500000 315.650000 ;
      RECT 1057.500000 314.350000 1058.500000 315.650000 ;
      RECT 1016.500000 314.350000 1049.500000 315.650000 ;
      RECT 1007.500000 314.350000 1008.500000 315.650000 ;
      RECT 966.500000 314.350000 999.500000 315.650000 ;
      RECT 957.500000 314.350000 958.500000 315.650000 ;
      RECT 916.500000 314.350000 949.500000 315.650000 ;
      RECT 907.500000 314.350000 908.500000 315.650000 ;
      RECT 866.500000 314.350000 899.500000 315.650000 ;
      RECT 857.500000 314.350000 858.500000 315.650000 ;
      RECT 816.500000 314.350000 849.500000 315.650000 ;
      RECT 807.500000 314.350000 808.500000 315.650000 ;
      RECT 766.500000 314.350000 799.500000 315.650000 ;
      RECT 757.500000 314.350000 758.500000 315.650000 ;
      RECT 716.500000 314.350000 749.500000 315.650000 ;
      RECT 707.500000 314.350000 708.500000 315.650000 ;
      RECT 666.500000 314.350000 699.500000 315.650000 ;
      RECT 657.500000 314.350000 658.500000 315.650000 ;
      RECT 616.500000 314.350000 649.500000 315.650000 ;
      RECT 607.500000 314.350000 608.500000 315.650000 ;
      RECT 566.500000 314.350000 599.500000 315.650000 ;
      RECT 557.500000 314.350000 558.500000 315.650000 ;
      RECT 516.500000 314.350000 549.500000 315.650000 ;
      RECT 507.500000 314.350000 508.500000 315.650000 ;
      RECT 416.500000 314.350000 499.500000 315.650000 ;
      RECT 407.500000 314.350000 408.500000 315.650000 ;
      RECT 366.500000 314.350000 399.500000 315.650000 ;
      RECT 357.500000 314.350000 358.500000 315.650000 ;
      RECT 316.500000 314.350000 349.500000 315.650000 ;
      RECT 307.500000 314.350000 308.500000 315.650000 ;
      RECT 266.500000 314.350000 299.500000 315.650000 ;
      RECT 257.500000 314.350000 258.500000 315.650000 ;
      RECT 216.500000 314.350000 249.500000 315.650000 ;
      RECT 207.500000 314.350000 208.500000 315.650000 ;
      RECT 166.500000 314.350000 199.500000 315.650000 ;
      RECT 157.500000 314.350000 158.500000 315.650000 ;
      RECT 116.500000 314.350000 149.500000 315.650000 ;
      RECT 107.500000 314.350000 108.500000 315.650000 ;
      RECT 66.500000 314.350000 99.500000 315.650000 ;
      RECT 57.500000 314.350000 58.500000 315.650000 ;
      RECT 29.500000 314.350000 49.500000 315.650000 ;
      RECT 15.500000 314.350000 16.500000 315.650000 ;
      RECT 1157.500000 313.650000 1170.500000 314.350000 ;
      RECT 1107.500000 313.650000 1149.500000 314.350000 ;
      RECT 1057.500000 313.650000 1099.500000 314.350000 ;
      RECT 1007.500000 313.650000 1049.500000 314.350000 ;
      RECT 957.500000 313.650000 999.500000 314.350000 ;
      RECT 907.500000 313.650000 949.500000 314.350000 ;
      RECT 857.500000 313.650000 899.500000 314.350000 ;
      RECT 807.500000 313.650000 849.500000 314.350000 ;
      RECT 757.500000 313.650000 799.500000 314.350000 ;
      RECT 707.500000 313.650000 749.500000 314.350000 ;
      RECT 657.500000 313.650000 699.500000 314.350000 ;
      RECT 607.500000 313.650000 649.500000 314.350000 ;
      RECT 557.500000 313.650000 599.500000 314.350000 ;
      RECT 507.500000 313.650000 549.500000 314.350000 ;
      RECT 407.500000 313.650000 499.500000 314.350000 ;
      RECT 357.500000 313.650000 399.500000 314.350000 ;
      RECT 307.500000 313.650000 349.500000 314.350000 ;
      RECT 257.500000 313.650000 299.500000 314.350000 ;
      RECT 207.500000 313.650000 249.500000 314.350000 ;
      RECT 157.500000 313.650000 199.500000 314.350000 ;
      RECT 107.500000 313.650000 149.500000 314.350000 ;
      RECT 57.500000 313.650000 99.500000 314.350000 ;
      RECT 15.500000 313.650000 49.500000 314.350000 ;
      RECT 1183.500000 312.350000 1186.000000 315.650000 ;
      RECT 1169.500000 312.350000 1170.500000 313.650000 ;
      RECT 1116.500000 312.350000 1149.500000 313.650000 ;
      RECT 1107.500000 312.350000 1108.500000 313.650000 ;
      RECT 1066.500000 312.350000 1099.500000 313.650000 ;
      RECT 1057.500000 312.350000 1058.500000 313.650000 ;
      RECT 1016.500000 312.350000 1049.500000 313.650000 ;
      RECT 1007.500000 312.350000 1008.500000 313.650000 ;
      RECT 966.500000 312.350000 999.500000 313.650000 ;
      RECT 957.500000 312.350000 958.500000 313.650000 ;
      RECT 916.500000 312.350000 949.500000 313.650000 ;
      RECT 907.500000 312.350000 908.500000 313.650000 ;
      RECT 866.500000 312.350000 899.500000 313.650000 ;
      RECT 857.500000 312.350000 858.500000 313.650000 ;
      RECT 816.500000 312.350000 849.500000 313.650000 ;
      RECT 807.500000 312.350000 808.500000 313.650000 ;
      RECT 766.500000 312.350000 799.500000 313.650000 ;
      RECT 757.500000 312.350000 758.500000 313.650000 ;
      RECT 716.500000 312.350000 749.500000 313.650000 ;
      RECT 707.500000 312.350000 708.500000 313.650000 ;
      RECT 666.500000 312.350000 699.500000 313.650000 ;
      RECT 657.500000 312.350000 658.500000 313.650000 ;
      RECT 616.500000 312.350000 649.500000 313.650000 ;
      RECT 607.500000 312.350000 608.500000 313.650000 ;
      RECT 566.500000 312.350000 599.500000 313.650000 ;
      RECT 557.500000 312.350000 558.500000 313.650000 ;
      RECT 516.500000 312.350000 549.500000 313.650000 ;
      RECT 507.500000 312.350000 508.500000 313.650000 ;
      RECT 416.500000 312.350000 499.500000 313.650000 ;
      RECT 407.500000 312.350000 408.500000 313.650000 ;
      RECT 366.500000 312.350000 399.500000 313.650000 ;
      RECT 357.500000 312.350000 358.500000 313.650000 ;
      RECT 316.500000 312.350000 349.500000 313.650000 ;
      RECT 307.500000 312.350000 308.500000 313.650000 ;
      RECT 266.500000 312.350000 299.500000 313.650000 ;
      RECT 257.500000 312.350000 258.500000 313.650000 ;
      RECT 216.500000 312.350000 249.500000 313.650000 ;
      RECT 207.500000 312.350000 208.500000 313.650000 ;
      RECT 166.500000 312.350000 199.500000 313.650000 ;
      RECT 157.500000 312.350000 158.500000 313.650000 ;
      RECT 116.500000 312.350000 149.500000 313.650000 ;
      RECT 107.500000 312.350000 108.500000 313.650000 ;
      RECT 66.500000 312.350000 99.500000 313.650000 ;
      RECT 57.500000 312.350000 58.500000 313.650000 ;
      RECT 29.500000 312.350000 49.500000 313.650000 ;
      RECT 15.500000 312.350000 16.500000 313.650000 ;
      RECT 0.000000 312.350000 2.500000 315.650000 ;
      RECT 1169.500000 311.650000 1186.000000 312.350000 ;
      RECT 1116.500000 311.650000 1156.500000 312.350000 ;
      RECT 1066.500000 311.650000 1108.500000 312.350000 ;
      RECT 1016.500000 311.650000 1058.500000 312.350000 ;
      RECT 966.500000 311.650000 1008.500000 312.350000 ;
      RECT 916.500000 311.650000 958.500000 312.350000 ;
      RECT 866.500000 311.650000 908.500000 312.350000 ;
      RECT 816.500000 311.650000 858.500000 312.350000 ;
      RECT 766.500000 311.650000 808.500000 312.350000 ;
      RECT 716.500000 311.650000 758.500000 312.350000 ;
      RECT 666.500000 311.650000 708.500000 312.350000 ;
      RECT 616.500000 311.650000 658.500000 312.350000 ;
      RECT 566.500000 311.650000 608.500000 312.350000 ;
      RECT 516.500000 311.650000 558.500000 312.350000 ;
      RECT 416.500000 311.650000 508.500000 312.350000 ;
      RECT 366.500000 311.650000 408.500000 312.350000 ;
      RECT 316.500000 311.650000 358.500000 312.350000 ;
      RECT 266.500000 311.650000 308.500000 312.350000 ;
      RECT 216.500000 311.650000 258.500000 312.350000 ;
      RECT 166.500000 311.650000 208.500000 312.350000 ;
      RECT 116.500000 311.650000 158.500000 312.350000 ;
      RECT 66.500000 311.650000 108.500000 312.350000 ;
      RECT 29.500000 311.650000 58.500000 312.350000 ;
      RECT 0.000000 311.650000 16.500000 312.350000 ;
      RECT 0.000000 311.170000 2.500000 311.650000 ;
      RECT 1183.500000 311.165000 1186.000000 311.650000 ;
      RECT 1169.500000 310.350000 1170.500000 311.650000 ;
      RECT 1116.500000 310.350000 1149.500000 311.650000 ;
      RECT 1107.500000 310.350000 1108.500000 311.650000 ;
      RECT 1066.500000 310.350000 1099.500000 311.650000 ;
      RECT 1057.500000 310.350000 1058.500000 311.650000 ;
      RECT 1016.500000 310.350000 1049.500000 311.650000 ;
      RECT 1007.500000 310.350000 1008.500000 311.650000 ;
      RECT 966.500000 310.350000 999.500000 311.650000 ;
      RECT 957.500000 310.350000 958.500000 311.650000 ;
      RECT 916.500000 310.350000 949.500000 311.650000 ;
      RECT 907.500000 310.350000 908.500000 311.650000 ;
      RECT 866.500000 310.350000 899.500000 311.650000 ;
      RECT 857.500000 310.350000 858.500000 311.650000 ;
      RECT 816.500000 310.350000 849.500000 311.650000 ;
      RECT 807.500000 310.350000 808.500000 311.650000 ;
      RECT 766.500000 310.350000 799.500000 311.650000 ;
      RECT 757.500000 310.350000 758.500000 311.650000 ;
      RECT 716.500000 310.350000 749.500000 311.650000 ;
      RECT 707.500000 310.350000 708.500000 311.650000 ;
      RECT 666.500000 310.350000 699.500000 311.650000 ;
      RECT 657.500000 310.350000 658.500000 311.650000 ;
      RECT 616.500000 310.350000 649.500000 311.650000 ;
      RECT 607.500000 310.350000 608.500000 311.650000 ;
      RECT 566.500000 310.350000 599.500000 311.650000 ;
      RECT 557.500000 310.350000 558.500000 311.650000 ;
      RECT 516.500000 310.350000 549.500000 311.650000 ;
      RECT 507.500000 310.350000 508.500000 311.650000 ;
      RECT 416.500000 310.350000 499.500000 311.650000 ;
      RECT 407.500000 310.350000 408.500000 311.650000 ;
      RECT 366.500000 310.350000 399.500000 311.650000 ;
      RECT 357.500000 310.350000 358.500000 311.650000 ;
      RECT 316.500000 310.350000 349.500000 311.650000 ;
      RECT 307.500000 310.350000 308.500000 311.650000 ;
      RECT 266.500000 310.350000 299.500000 311.650000 ;
      RECT 257.500000 310.350000 258.500000 311.650000 ;
      RECT 216.500000 310.350000 249.500000 311.650000 ;
      RECT 207.500000 310.350000 208.500000 311.650000 ;
      RECT 166.500000 310.350000 199.500000 311.650000 ;
      RECT 157.500000 310.350000 158.500000 311.650000 ;
      RECT 116.500000 310.350000 149.500000 311.650000 ;
      RECT 107.500000 310.350000 108.500000 311.650000 ;
      RECT 66.500000 310.350000 99.500000 311.650000 ;
      RECT 57.500000 310.350000 58.500000 311.650000 ;
      RECT 29.500000 310.350000 49.500000 311.650000 ;
      RECT 15.500000 310.350000 16.500000 311.650000 ;
      RECT 1157.500000 309.650000 1170.500000 310.350000 ;
      RECT 1107.500000 309.650000 1149.500000 310.350000 ;
      RECT 1057.500000 309.650000 1099.500000 310.350000 ;
      RECT 1007.500000 309.650000 1049.500000 310.350000 ;
      RECT 957.500000 309.650000 999.500000 310.350000 ;
      RECT 907.500000 309.650000 949.500000 310.350000 ;
      RECT 857.500000 309.650000 899.500000 310.350000 ;
      RECT 807.500000 309.650000 849.500000 310.350000 ;
      RECT 757.500000 309.650000 799.500000 310.350000 ;
      RECT 707.500000 309.650000 749.500000 310.350000 ;
      RECT 657.500000 309.650000 699.500000 310.350000 ;
      RECT 607.500000 309.650000 649.500000 310.350000 ;
      RECT 557.500000 309.650000 599.500000 310.350000 ;
      RECT 507.500000 309.650000 549.500000 310.350000 ;
      RECT 407.500000 309.650000 499.500000 310.350000 ;
      RECT 357.500000 309.650000 399.500000 310.350000 ;
      RECT 307.500000 309.650000 349.500000 310.350000 ;
      RECT 257.500000 309.650000 299.500000 310.350000 ;
      RECT 207.500000 309.650000 249.500000 310.350000 ;
      RECT 157.500000 309.650000 199.500000 310.350000 ;
      RECT 107.500000 309.650000 149.500000 310.350000 ;
      RECT 57.500000 309.650000 99.500000 310.350000 ;
      RECT 15.500000 309.650000 49.500000 310.350000 ;
      RECT 1183.500000 308.350000 1183.980000 311.165000 ;
      RECT 1169.500000 308.350000 1170.500000 309.650000 ;
      RECT 1116.500000 308.350000 1149.500000 309.650000 ;
      RECT 1107.500000 308.350000 1108.500000 309.650000 ;
      RECT 1066.500000 308.350000 1099.500000 309.650000 ;
      RECT 1057.500000 308.350000 1058.500000 309.650000 ;
      RECT 1016.500000 308.350000 1049.500000 309.650000 ;
      RECT 1007.500000 308.350000 1008.500000 309.650000 ;
      RECT 966.500000 308.350000 999.500000 309.650000 ;
      RECT 957.500000 308.350000 958.500000 309.650000 ;
      RECT 916.500000 308.350000 949.500000 309.650000 ;
      RECT 907.500000 308.350000 908.500000 309.650000 ;
      RECT 866.500000 308.350000 899.500000 309.650000 ;
      RECT 857.500000 308.350000 858.500000 309.650000 ;
      RECT 816.500000 308.350000 849.500000 309.650000 ;
      RECT 807.500000 308.350000 808.500000 309.650000 ;
      RECT 766.500000 308.350000 799.500000 309.650000 ;
      RECT 757.500000 308.350000 758.500000 309.650000 ;
      RECT 716.500000 308.350000 749.500000 309.650000 ;
      RECT 707.500000 308.350000 708.500000 309.650000 ;
      RECT 666.500000 308.350000 699.500000 309.650000 ;
      RECT 657.500000 308.350000 658.500000 309.650000 ;
      RECT 616.500000 308.350000 649.500000 309.650000 ;
      RECT 607.500000 308.350000 608.500000 309.650000 ;
      RECT 566.500000 308.350000 599.500000 309.650000 ;
      RECT 557.500000 308.350000 558.500000 309.650000 ;
      RECT 516.500000 308.350000 549.500000 309.650000 ;
      RECT 507.500000 308.350000 508.500000 309.650000 ;
      RECT 416.500000 308.350000 499.500000 309.650000 ;
      RECT 407.500000 308.350000 408.500000 309.650000 ;
      RECT 366.500000 308.350000 399.500000 309.650000 ;
      RECT 357.500000 308.350000 358.500000 309.650000 ;
      RECT 316.500000 308.350000 349.500000 309.650000 ;
      RECT 307.500000 308.350000 308.500000 309.650000 ;
      RECT 266.500000 308.350000 299.500000 309.650000 ;
      RECT 257.500000 308.350000 258.500000 309.650000 ;
      RECT 216.500000 308.350000 249.500000 309.650000 ;
      RECT 207.500000 308.350000 208.500000 309.650000 ;
      RECT 166.500000 308.350000 199.500000 309.650000 ;
      RECT 157.500000 308.350000 158.500000 309.650000 ;
      RECT 116.500000 308.350000 149.500000 309.650000 ;
      RECT 107.500000 308.350000 108.500000 309.650000 ;
      RECT 66.500000 308.350000 99.500000 309.650000 ;
      RECT 57.500000 308.350000 58.500000 309.650000 ;
      RECT 29.500000 308.350000 49.500000 309.650000 ;
      RECT 15.500000 308.350000 16.500000 309.650000 ;
      RECT 2.020000 308.350000 2.500000 311.170000 ;
      RECT 2.020000 308.070000 16.500000 308.350000 ;
      RECT 1169.500000 308.065000 1183.980000 308.350000 ;
      RECT 1169.500000 307.650000 1186.000000 308.065000 ;
      RECT 1116.500000 307.650000 1156.500000 308.350000 ;
      RECT 1066.500000 307.650000 1108.500000 308.350000 ;
      RECT 1016.500000 307.650000 1058.500000 308.350000 ;
      RECT 966.500000 307.650000 1008.500000 308.350000 ;
      RECT 916.500000 307.650000 958.500000 308.350000 ;
      RECT 866.500000 307.650000 908.500000 308.350000 ;
      RECT 816.500000 307.650000 858.500000 308.350000 ;
      RECT 766.500000 307.650000 808.500000 308.350000 ;
      RECT 716.500000 307.650000 758.500000 308.350000 ;
      RECT 666.500000 307.650000 708.500000 308.350000 ;
      RECT 616.500000 307.650000 658.500000 308.350000 ;
      RECT 566.500000 307.650000 608.500000 308.350000 ;
      RECT 516.500000 307.650000 558.500000 308.350000 ;
      RECT 416.500000 307.650000 508.500000 308.350000 ;
      RECT 366.500000 307.650000 408.500000 308.350000 ;
      RECT 316.500000 307.650000 358.500000 308.350000 ;
      RECT 266.500000 307.650000 308.500000 308.350000 ;
      RECT 216.500000 307.650000 258.500000 308.350000 ;
      RECT 166.500000 307.650000 208.500000 308.350000 ;
      RECT 116.500000 307.650000 158.500000 308.350000 ;
      RECT 66.500000 307.650000 108.500000 308.350000 ;
      RECT 29.500000 307.650000 58.500000 308.350000 ;
      RECT 0.000000 307.650000 16.500000 308.070000 ;
      RECT 1169.500000 306.350000 1170.500000 307.650000 ;
      RECT 1116.500000 306.350000 1149.500000 307.650000 ;
      RECT 1107.500000 306.350000 1108.500000 307.650000 ;
      RECT 1066.500000 306.350000 1099.500000 307.650000 ;
      RECT 1057.500000 306.350000 1058.500000 307.650000 ;
      RECT 1016.500000 306.350000 1049.500000 307.650000 ;
      RECT 1007.500000 306.350000 1008.500000 307.650000 ;
      RECT 966.500000 306.350000 999.500000 307.650000 ;
      RECT 957.500000 306.350000 958.500000 307.650000 ;
      RECT 916.500000 306.350000 949.500000 307.650000 ;
      RECT 907.500000 306.350000 908.500000 307.650000 ;
      RECT 866.500000 306.350000 899.500000 307.650000 ;
      RECT 857.500000 306.350000 858.500000 307.650000 ;
      RECT 816.500000 306.350000 849.500000 307.650000 ;
      RECT 807.500000 306.350000 808.500000 307.650000 ;
      RECT 766.500000 306.350000 799.500000 307.650000 ;
      RECT 757.500000 306.350000 758.500000 307.650000 ;
      RECT 716.500000 306.350000 749.500000 307.650000 ;
      RECT 707.500000 306.350000 708.500000 307.650000 ;
      RECT 666.500000 306.350000 699.500000 307.650000 ;
      RECT 657.500000 306.350000 658.500000 307.650000 ;
      RECT 616.500000 306.350000 649.500000 307.650000 ;
      RECT 607.500000 306.350000 608.500000 307.650000 ;
      RECT 566.500000 306.350000 599.500000 307.650000 ;
      RECT 557.500000 306.350000 558.500000 307.650000 ;
      RECT 516.500000 306.350000 549.500000 307.650000 ;
      RECT 507.500000 306.350000 508.500000 307.650000 ;
      RECT 416.500000 306.350000 499.500000 307.650000 ;
      RECT 407.500000 306.350000 408.500000 307.650000 ;
      RECT 366.500000 306.350000 399.500000 307.650000 ;
      RECT 357.500000 306.350000 358.500000 307.650000 ;
      RECT 316.500000 306.350000 349.500000 307.650000 ;
      RECT 307.500000 306.350000 308.500000 307.650000 ;
      RECT 266.500000 306.350000 299.500000 307.650000 ;
      RECT 257.500000 306.350000 258.500000 307.650000 ;
      RECT 216.500000 306.350000 249.500000 307.650000 ;
      RECT 207.500000 306.350000 208.500000 307.650000 ;
      RECT 166.500000 306.350000 199.500000 307.650000 ;
      RECT 157.500000 306.350000 158.500000 307.650000 ;
      RECT 116.500000 306.350000 149.500000 307.650000 ;
      RECT 107.500000 306.350000 108.500000 307.650000 ;
      RECT 66.500000 306.350000 99.500000 307.650000 ;
      RECT 57.500000 306.350000 58.500000 307.650000 ;
      RECT 29.500000 306.350000 49.500000 307.650000 ;
      RECT 15.500000 306.350000 16.500000 307.650000 ;
      RECT 1157.500000 305.650000 1170.500000 306.350000 ;
      RECT 1107.500000 305.650000 1149.500000 306.350000 ;
      RECT 1057.500000 305.650000 1099.500000 306.350000 ;
      RECT 1007.500000 305.650000 1049.500000 306.350000 ;
      RECT 957.500000 305.650000 999.500000 306.350000 ;
      RECT 907.500000 305.650000 949.500000 306.350000 ;
      RECT 857.500000 305.650000 899.500000 306.350000 ;
      RECT 807.500000 305.650000 849.500000 306.350000 ;
      RECT 757.500000 305.650000 799.500000 306.350000 ;
      RECT 707.500000 305.650000 749.500000 306.350000 ;
      RECT 657.500000 305.650000 699.500000 306.350000 ;
      RECT 607.500000 305.650000 649.500000 306.350000 ;
      RECT 557.500000 305.650000 599.500000 306.350000 ;
      RECT 507.500000 305.650000 549.500000 306.350000 ;
      RECT 407.500000 305.650000 499.500000 306.350000 ;
      RECT 357.500000 305.650000 399.500000 306.350000 ;
      RECT 307.500000 305.650000 349.500000 306.350000 ;
      RECT 257.500000 305.650000 299.500000 306.350000 ;
      RECT 207.500000 305.650000 249.500000 306.350000 ;
      RECT 157.500000 305.650000 199.500000 306.350000 ;
      RECT 107.500000 305.650000 149.500000 306.350000 ;
      RECT 57.500000 305.650000 99.500000 306.350000 ;
      RECT 15.500000 305.650000 49.500000 306.350000 ;
      RECT 1183.500000 305.485000 1186.000000 307.650000 ;
      RECT 1183.500000 304.350000 1183.980000 305.485000 ;
      RECT 1169.500000 304.350000 1170.500000 305.650000 ;
      RECT 1116.500000 304.350000 1149.500000 305.650000 ;
      RECT 1107.500000 304.350000 1108.500000 305.650000 ;
      RECT 1066.500000 304.350000 1099.500000 305.650000 ;
      RECT 1057.500000 304.350000 1058.500000 305.650000 ;
      RECT 1016.500000 304.350000 1049.500000 305.650000 ;
      RECT 1007.500000 304.350000 1008.500000 305.650000 ;
      RECT 966.500000 304.350000 999.500000 305.650000 ;
      RECT 957.500000 304.350000 958.500000 305.650000 ;
      RECT 916.500000 304.350000 949.500000 305.650000 ;
      RECT 907.500000 304.350000 908.500000 305.650000 ;
      RECT 866.500000 304.350000 899.500000 305.650000 ;
      RECT 857.500000 304.350000 858.500000 305.650000 ;
      RECT 816.500000 304.350000 849.500000 305.650000 ;
      RECT 807.500000 304.350000 808.500000 305.650000 ;
      RECT 766.500000 304.350000 799.500000 305.650000 ;
      RECT 757.500000 304.350000 758.500000 305.650000 ;
      RECT 716.500000 304.350000 749.500000 305.650000 ;
      RECT 707.500000 304.350000 708.500000 305.650000 ;
      RECT 666.500000 304.350000 699.500000 305.650000 ;
      RECT 657.500000 304.350000 658.500000 305.650000 ;
      RECT 616.500000 304.350000 649.500000 305.650000 ;
      RECT 607.500000 304.350000 608.500000 305.650000 ;
      RECT 566.500000 304.350000 599.500000 305.650000 ;
      RECT 557.500000 304.350000 558.500000 305.650000 ;
      RECT 516.500000 304.350000 549.500000 305.650000 ;
      RECT 507.500000 304.350000 508.500000 305.650000 ;
      RECT 416.500000 304.350000 499.500000 305.650000 ;
      RECT 407.500000 304.350000 408.500000 305.650000 ;
      RECT 366.500000 304.350000 399.500000 305.650000 ;
      RECT 357.500000 304.350000 358.500000 305.650000 ;
      RECT 316.500000 304.350000 349.500000 305.650000 ;
      RECT 307.500000 304.350000 308.500000 305.650000 ;
      RECT 266.500000 304.350000 299.500000 305.650000 ;
      RECT 257.500000 304.350000 258.500000 305.650000 ;
      RECT 216.500000 304.350000 249.500000 305.650000 ;
      RECT 207.500000 304.350000 208.500000 305.650000 ;
      RECT 166.500000 304.350000 199.500000 305.650000 ;
      RECT 157.500000 304.350000 158.500000 305.650000 ;
      RECT 116.500000 304.350000 149.500000 305.650000 ;
      RECT 107.500000 304.350000 108.500000 305.650000 ;
      RECT 66.500000 304.350000 99.500000 305.650000 ;
      RECT 57.500000 304.350000 58.500000 305.650000 ;
      RECT 29.500000 304.350000 49.500000 305.650000 ;
      RECT 15.500000 304.350000 16.500000 305.650000 ;
      RECT 0.000000 304.350000 2.500000 307.650000 ;
      RECT 1169.500000 303.650000 1183.980000 304.350000 ;
      RECT 1116.500000 303.650000 1156.500000 304.350000 ;
      RECT 1066.500000 303.650000 1108.500000 304.350000 ;
      RECT 1016.500000 303.650000 1058.500000 304.350000 ;
      RECT 966.500000 303.650000 1008.500000 304.350000 ;
      RECT 916.500000 303.650000 958.500000 304.350000 ;
      RECT 866.500000 303.650000 908.500000 304.350000 ;
      RECT 816.500000 303.650000 858.500000 304.350000 ;
      RECT 766.500000 303.650000 808.500000 304.350000 ;
      RECT 716.500000 303.650000 758.500000 304.350000 ;
      RECT 666.500000 303.650000 708.500000 304.350000 ;
      RECT 616.500000 303.650000 658.500000 304.350000 ;
      RECT 566.500000 303.650000 608.500000 304.350000 ;
      RECT 516.500000 303.650000 558.500000 304.350000 ;
      RECT 416.500000 303.650000 508.500000 304.350000 ;
      RECT 366.500000 303.650000 408.500000 304.350000 ;
      RECT 316.500000 303.650000 358.500000 304.350000 ;
      RECT 266.500000 303.650000 308.500000 304.350000 ;
      RECT 216.500000 303.650000 258.500000 304.350000 ;
      RECT 166.500000 303.650000 208.500000 304.350000 ;
      RECT 116.500000 303.650000 158.500000 304.350000 ;
      RECT 66.500000 303.650000 108.500000 304.350000 ;
      RECT 29.500000 303.650000 58.500000 304.350000 ;
      RECT 0.000000 303.650000 16.500000 304.350000 ;
      RECT 1183.500000 302.385000 1183.980000 303.650000 ;
      RECT 1169.500000 302.350000 1170.500000 303.650000 ;
      RECT 1116.500000 302.350000 1149.500000 303.650000 ;
      RECT 1107.500000 302.350000 1108.500000 303.650000 ;
      RECT 1066.500000 302.350000 1099.500000 303.650000 ;
      RECT 1057.500000 302.350000 1058.500000 303.650000 ;
      RECT 1016.500000 302.350000 1049.500000 303.650000 ;
      RECT 1007.500000 302.350000 1008.500000 303.650000 ;
      RECT 966.500000 302.350000 999.500000 303.650000 ;
      RECT 957.500000 302.350000 958.500000 303.650000 ;
      RECT 916.500000 302.350000 949.500000 303.650000 ;
      RECT 907.500000 302.350000 908.500000 303.650000 ;
      RECT 866.500000 302.350000 899.500000 303.650000 ;
      RECT 857.500000 302.350000 858.500000 303.650000 ;
      RECT 816.500000 302.350000 849.500000 303.650000 ;
      RECT 807.500000 302.350000 808.500000 303.650000 ;
      RECT 766.500000 302.350000 799.500000 303.650000 ;
      RECT 757.500000 302.350000 758.500000 303.650000 ;
      RECT 716.500000 302.350000 749.500000 303.650000 ;
      RECT 707.500000 302.350000 708.500000 303.650000 ;
      RECT 666.500000 302.350000 699.500000 303.650000 ;
      RECT 657.500000 302.350000 658.500000 303.650000 ;
      RECT 616.500000 302.350000 649.500000 303.650000 ;
      RECT 607.500000 302.350000 608.500000 303.650000 ;
      RECT 566.500000 302.350000 599.500000 303.650000 ;
      RECT 557.500000 302.350000 558.500000 303.650000 ;
      RECT 516.500000 302.350000 549.500000 303.650000 ;
      RECT 507.500000 302.350000 508.500000 303.650000 ;
      RECT 416.500000 302.350000 499.500000 303.650000 ;
      RECT 407.500000 302.350000 408.500000 303.650000 ;
      RECT 366.500000 302.350000 399.500000 303.650000 ;
      RECT 357.500000 302.350000 358.500000 303.650000 ;
      RECT 316.500000 302.350000 349.500000 303.650000 ;
      RECT 307.500000 302.350000 308.500000 303.650000 ;
      RECT 266.500000 302.350000 299.500000 303.650000 ;
      RECT 257.500000 302.350000 258.500000 303.650000 ;
      RECT 216.500000 302.350000 249.500000 303.650000 ;
      RECT 207.500000 302.350000 208.500000 303.650000 ;
      RECT 166.500000 302.350000 199.500000 303.650000 ;
      RECT 157.500000 302.350000 158.500000 303.650000 ;
      RECT 116.500000 302.350000 149.500000 303.650000 ;
      RECT 107.500000 302.350000 108.500000 303.650000 ;
      RECT 66.500000 302.350000 99.500000 303.650000 ;
      RECT 57.500000 302.350000 58.500000 303.650000 ;
      RECT 29.500000 302.350000 49.500000 303.650000 ;
      RECT 15.500000 302.350000 16.500000 303.650000 ;
      RECT 1157.500000 301.650000 1170.500000 302.350000 ;
      RECT 1107.500000 301.650000 1149.500000 302.350000 ;
      RECT 1057.500000 301.650000 1099.500000 302.350000 ;
      RECT 1007.500000 301.650000 1049.500000 302.350000 ;
      RECT 957.500000 301.650000 999.500000 302.350000 ;
      RECT 907.500000 301.650000 949.500000 302.350000 ;
      RECT 857.500000 301.650000 899.500000 302.350000 ;
      RECT 807.500000 301.650000 849.500000 302.350000 ;
      RECT 757.500000 301.650000 799.500000 302.350000 ;
      RECT 707.500000 301.650000 749.500000 302.350000 ;
      RECT 657.500000 301.650000 699.500000 302.350000 ;
      RECT 607.500000 301.650000 649.500000 302.350000 ;
      RECT 557.500000 301.650000 599.500000 302.350000 ;
      RECT 507.500000 301.650000 549.500000 302.350000 ;
      RECT 407.500000 301.650000 499.500000 302.350000 ;
      RECT 357.500000 301.650000 399.500000 302.350000 ;
      RECT 307.500000 301.650000 349.500000 302.350000 ;
      RECT 257.500000 301.650000 299.500000 302.350000 ;
      RECT 207.500000 301.650000 249.500000 302.350000 ;
      RECT 157.500000 301.650000 199.500000 302.350000 ;
      RECT 107.500000 301.650000 149.500000 302.350000 ;
      RECT 57.500000 301.650000 99.500000 302.350000 ;
      RECT 15.500000 301.650000 49.500000 302.350000 ;
      RECT 1183.500000 301.525000 1186.000000 302.385000 ;
      RECT 0.000000 300.575000 2.500000 303.650000 ;
      RECT 1183.500000 300.350000 1183.980000 301.525000 ;
      RECT 1169.500000 300.350000 1170.500000 301.650000 ;
      RECT 1116.500000 300.350000 1149.500000 301.650000 ;
      RECT 1107.500000 300.350000 1108.500000 301.650000 ;
      RECT 1066.500000 300.350000 1099.500000 301.650000 ;
      RECT 1057.500000 300.350000 1058.500000 301.650000 ;
      RECT 1016.500000 300.350000 1049.500000 301.650000 ;
      RECT 1007.500000 300.350000 1008.500000 301.650000 ;
      RECT 966.500000 300.350000 999.500000 301.650000 ;
      RECT 957.500000 300.350000 958.500000 301.650000 ;
      RECT 916.500000 300.350000 949.500000 301.650000 ;
      RECT 907.500000 300.350000 908.500000 301.650000 ;
      RECT 866.500000 300.350000 899.500000 301.650000 ;
      RECT 857.500000 300.350000 858.500000 301.650000 ;
      RECT 816.500000 300.350000 849.500000 301.650000 ;
      RECT 807.500000 300.350000 808.500000 301.650000 ;
      RECT 766.500000 300.350000 799.500000 301.650000 ;
      RECT 757.500000 300.350000 758.500000 301.650000 ;
      RECT 716.500000 300.350000 749.500000 301.650000 ;
      RECT 707.500000 300.350000 708.500000 301.650000 ;
      RECT 666.500000 300.350000 699.500000 301.650000 ;
      RECT 657.500000 300.350000 658.500000 301.650000 ;
      RECT 616.500000 300.350000 649.500000 301.650000 ;
      RECT 607.500000 300.350000 608.500000 301.650000 ;
      RECT 566.500000 300.350000 599.500000 301.650000 ;
      RECT 557.500000 300.350000 558.500000 301.650000 ;
      RECT 516.500000 300.350000 549.500000 301.650000 ;
      RECT 507.500000 300.350000 508.500000 301.650000 ;
      RECT 416.500000 300.350000 499.500000 301.650000 ;
      RECT 407.500000 300.350000 408.500000 301.650000 ;
      RECT 366.500000 300.350000 399.500000 301.650000 ;
      RECT 357.500000 300.350000 358.500000 301.650000 ;
      RECT 316.500000 300.350000 349.500000 301.650000 ;
      RECT 307.500000 300.350000 308.500000 301.650000 ;
      RECT 266.500000 300.350000 299.500000 301.650000 ;
      RECT 257.500000 300.350000 258.500000 301.650000 ;
      RECT 216.500000 300.350000 249.500000 301.650000 ;
      RECT 207.500000 300.350000 208.500000 301.650000 ;
      RECT 166.500000 300.350000 199.500000 301.650000 ;
      RECT 157.500000 300.350000 158.500000 301.650000 ;
      RECT 116.500000 300.350000 149.500000 301.650000 ;
      RECT 107.500000 300.350000 108.500000 301.650000 ;
      RECT 66.500000 300.350000 99.500000 301.650000 ;
      RECT 57.500000 300.350000 58.500000 301.650000 ;
      RECT 29.500000 300.350000 49.500000 301.650000 ;
      RECT 15.500000 300.350000 16.500000 301.650000 ;
      RECT 2.020000 300.350000 2.500000 300.575000 ;
      RECT 1169.500000 299.650000 1183.980000 300.350000 ;
      RECT 1116.500000 299.650000 1156.500000 300.350000 ;
      RECT 1066.500000 299.650000 1108.500000 300.350000 ;
      RECT 1016.500000 299.650000 1058.500000 300.350000 ;
      RECT 966.500000 299.650000 1008.500000 300.350000 ;
      RECT 916.500000 299.650000 958.500000 300.350000 ;
      RECT 866.500000 299.650000 908.500000 300.350000 ;
      RECT 816.500000 299.650000 858.500000 300.350000 ;
      RECT 766.500000 299.650000 808.500000 300.350000 ;
      RECT 716.500000 299.650000 758.500000 300.350000 ;
      RECT 666.500000 299.650000 708.500000 300.350000 ;
      RECT 616.500000 299.650000 658.500000 300.350000 ;
      RECT 566.500000 299.650000 608.500000 300.350000 ;
      RECT 516.500000 299.650000 558.500000 300.350000 ;
      RECT 416.500000 299.650000 508.500000 300.350000 ;
      RECT 366.500000 299.650000 408.500000 300.350000 ;
      RECT 316.500000 299.650000 358.500000 300.350000 ;
      RECT 266.500000 299.650000 308.500000 300.350000 ;
      RECT 216.500000 299.650000 258.500000 300.350000 ;
      RECT 166.500000 299.650000 208.500000 300.350000 ;
      RECT 116.500000 299.650000 158.500000 300.350000 ;
      RECT 66.500000 299.650000 108.500000 300.350000 ;
      RECT 29.500000 299.650000 58.500000 300.350000 ;
      RECT 2.020000 299.650000 16.500000 300.350000 ;
      RECT 1183.500000 298.425000 1183.980000 299.650000 ;
      RECT 1169.500000 298.350000 1170.500000 299.650000 ;
      RECT 1116.500000 298.350000 1149.500000 299.650000 ;
      RECT 1107.500000 298.350000 1108.500000 299.650000 ;
      RECT 1066.500000 298.350000 1099.500000 299.650000 ;
      RECT 1057.500000 298.350000 1058.500000 299.650000 ;
      RECT 1016.500000 298.350000 1049.500000 299.650000 ;
      RECT 1007.500000 298.350000 1008.500000 299.650000 ;
      RECT 966.500000 298.350000 999.500000 299.650000 ;
      RECT 957.500000 298.350000 958.500000 299.650000 ;
      RECT 916.500000 298.350000 949.500000 299.650000 ;
      RECT 907.500000 298.350000 908.500000 299.650000 ;
      RECT 866.500000 298.350000 899.500000 299.650000 ;
      RECT 857.500000 298.350000 858.500000 299.650000 ;
      RECT 816.500000 298.350000 849.500000 299.650000 ;
      RECT 807.500000 298.350000 808.500000 299.650000 ;
      RECT 766.500000 298.350000 799.500000 299.650000 ;
      RECT 757.500000 298.350000 758.500000 299.650000 ;
      RECT 716.500000 298.350000 749.500000 299.650000 ;
      RECT 707.500000 298.350000 708.500000 299.650000 ;
      RECT 666.500000 298.350000 699.500000 299.650000 ;
      RECT 657.500000 298.350000 658.500000 299.650000 ;
      RECT 616.500000 298.350000 649.500000 299.650000 ;
      RECT 607.500000 298.350000 608.500000 299.650000 ;
      RECT 566.500000 298.350000 599.500000 299.650000 ;
      RECT 557.500000 298.350000 558.500000 299.650000 ;
      RECT 516.500000 298.350000 549.500000 299.650000 ;
      RECT 507.500000 298.350000 508.500000 299.650000 ;
      RECT 416.500000 298.350000 449.500000 299.650000 ;
      RECT 407.500000 298.350000 408.500000 299.650000 ;
      RECT 366.500000 298.350000 399.500000 299.650000 ;
      RECT 357.500000 298.350000 358.500000 299.650000 ;
      RECT 316.500000 298.350000 349.500000 299.650000 ;
      RECT 307.500000 298.350000 308.500000 299.650000 ;
      RECT 266.500000 298.350000 299.500000 299.650000 ;
      RECT 257.500000 298.350000 258.500000 299.650000 ;
      RECT 216.500000 298.350000 249.500000 299.650000 ;
      RECT 207.500000 298.350000 208.500000 299.650000 ;
      RECT 166.500000 298.350000 199.500000 299.650000 ;
      RECT 157.500000 298.350000 158.500000 299.650000 ;
      RECT 116.500000 298.350000 149.500000 299.650000 ;
      RECT 107.500000 298.350000 108.500000 299.650000 ;
      RECT 66.500000 298.350000 99.500000 299.650000 ;
      RECT 57.500000 298.350000 58.500000 299.650000 ;
      RECT 29.500000 298.350000 49.500000 299.650000 ;
      RECT 15.500000 298.350000 16.500000 299.650000 ;
      RECT 1157.500000 297.650000 1170.500000 298.350000 ;
      RECT 1107.500000 297.650000 1149.500000 298.350000 ;
      RECT 1057.500000 297.650000 1099.500000 298.350000 ;
      RECT 1007.500000 297.650000 1049.500000 298.350000 ;
      RECT 957.500000 297.650000 999.500000 298.350000 ;
      RECT 907.500000 297.650000 949.500000 298.350000 ;
      RECT 857.500000 297.650000 899.500000 298.350000 ;
      RECT 807.500000 297.650000 849.500000 298.350000 ;
      RECT 757.500000 297.650000 799.500000 298.350000 ;
      RECT 707.500000 297.650000 749.500000 298.350000 ;
      RECT 657.500000 297.650000 699.500000 298.350000 ;
      RECT 607.500000 297.650000 649.500000 298.350000 ;
      RECT 557.500000 297.650000 599.500000 298.350000 ;
      RECT 507.500000 297.650000 549.500000 298.350000 ;
      RECT 457.500000 297.650000 499.500000 299.650000 ;
      RECT 407.500000 297.650000 449.500000 298.350000 ;
      RECT 357.500000 297.650000 399.500000 298.350000 ;
      RECT 307.500000 297.650000 349.500000 298.350000 ;
      RECT 257.500000 297.650000 299.500000 298.350000 ;
      RECT 207.500000 297.650000 249.500000 298.350000 ;
      RECT 157.500000 297.650000 199.500000 298.350000 ;
      RECT 107.500000 297.650000 149.500000 298.350000 ;
      RECT 57.500000 297.650000 99.500000 298.350000 ;
      RECT 15.500000 297.650000 49.500000 298.350000 ;
      RECT 2.020000 297.475000 2.500000 299.650000 ;
      RECT 0.000000 296.615000 2.500000 297.475000 ;
      RECT 1183.500000 296.350000 1186.000000 298.425000 ;
      RECT 1169.500000 296.350000 1170.500000 297.650000 ;
      RECT 1116.500000 296.350000 1149.500000 297.650000 ;
      RECT 1107.500000 296.350000 1108.500000 297.650000 ;
      RECT 1066.500000 296.350000 1099.500000 297.650000 ;
      RECT 1057.500000 296.350000 1058.500000 297.650000 ;
      RECT 1016.500000 296.350000 1049.500000 297.650000 ;
      RECT 1007.500000 296.350000 1008.500000 297.650000 ;
      RECT 966.500000 296.350000 999.500000 297.650000 ;
      RECT 957.500000 296.350000 958.500000 297.650000 ;
      RECT 916.500000 296.350000 949.500000 297.650000 ;
      RECT 907.500000 296.350000 908.500000 297.650000 ;
      RECT 866.500000 296.350000 899.500000 297.650000 ;
      RECT 857.500000 296.350000 858.500000 297.650000 ;
      RECT 816.500000 296.350000 849.500000 297.650000 ;
      RECT 807.500000 296.350000 808.500000 297.650000 ;
      RECT 766.500000 296.350000 799.500000 297.650000 ;
      RECT 757.500000 296.350000 758.500000 297.650000 ;
      RECT 716.500000 296.350000 749.500000 297.650000 ;
      RECT 707.500000 296.350000 708.500000 297.650000 ;
      RECT 666.500000 296.350000 699.500000 297.650000 ;
      RECT 657.500000 296.350000 658.500000 297.650000 ;
      RECT 616.500000 296.350000 649.500000 297.650000 ;
      RECT 607.500000 296.350000 608.500000 297.650000 ;
      RECT 566.500000 296.350000 599.500000 297.650000 ;
      RECT 557.500000 296.350000 558.500000 297.650000 ;
      RECT 516.500000 296.350000 549.500000 297.650000 ;
      RECT 507.500000 296.350000 508.500000 297.650000 ;
      RECT 466.500000 296.350000 499.500000 297.650000 ;
      RECT 457.500000 296.350000 458.500000 297.650000 ;
      RECT 416.500000 296.350000 449.500000 297.650000 ;
      RECT 407.500000 296.350000 408.500000 297.650000 ;
      RECT 366.500000 296.350000 399.500000 297.650000 ;
      RECT 357.500000 296.350000 358.500000 297.650000 ;
      RECT 316.500000 296.350000 349.500000 297.650000 ;
      RECT 307.500000 296.350000 308.500000 297.650000 ;
      RECT 266.500000 296.350000 299.500000 297.650000 ;
      RECT 257.500000 296.350000 258.500000 297.650000 ;
      RECT 216.500000 296.350000 249.500000 297.650000 ;
      RECT 207.500000 296.350000 208.500000 297.650000 ;
      RECT 166.500000 296.350000 199.500000 297.650000 ;
      RECT 157.500000 296.350000 158.500000 297.650000 ;
      RECT 116.500000 296.350000 149.500000 297.650000 ;
      RECT 107.500000 296.350000 108.500000 297.650000 ;
      RECT 66.500000 296.350000 99.500000 297.650000 ;
      RECT 57.500000 296.350000 58.500000 297.650000 ;
      RECT 29.500000 296.350000 49.500000 297.650000 ;
      RECT 15.500000 296.350000 16.500000 297.650000 ;
      RECT 2.020000 296.350000 2.500000 296.615000 ;
      RECT 1169.500000 295.650000 1186.000000 296.350000 ;
      RECT 1116.500000 295.650000 1156.500000 296.350000 ;
      RECT 1066.500000 295.650000 1108.500000 296.350000 ;
      RECT 1016.500000 295.650000 1058.500000 296.350000 ;
      RECT 966.500000 295.650000 1008.500000 296.350000 ;
      RECT 916.500000 295.650000 958.500000 296.350000 ;
      RECT 866.500000 295.650000 908.500000 296.350000 ;
      RECT 816.500000 295.650000 858.500000 296.350000 ;
      RECT 766.500000 295.650000 808.500000 296.350000 ;
      RECT 716.500000 295.650000 758.500000 296.350000 ;
      RECT 666.500000 295.650000 708.500000 296.350000 ;
      RECT 616.500000 295.650000 658.500000 296.350000 ;
      RECT 566.500000 295.650000 608.500000 296.350000 ;
      RECT 516.500000 295.650000 558.500000 296.350000 ;
      RECT 466.500000 295.650000 508.500000 296.350000 ;
      RECT 416.500000 295.650000 458.500000 296.350000 ;
      RECT 366.500000 295.650000 408.500000 296.350000 ;
      RECT 316.500000 295.650000 358.500000 296.350000 ;
      RECT 266.500000 295.650000 308.500000 296.350000 ;
      RECT 216.500000 295.650000 258.500000 296.350000 ;
      RECT 166.500000 295.650000 208.500000 296.350000 ;
      RECT 116.500000 295.650000 158.500000 296.350000 ;
      RECT 66.500000 295.650000 108.500000 296.350000 ;
      RECT 29.500000 295.650000 58.500000 296.350000 ;
      RECT 2.020000 295.650000 16.500000 296.350000 ;
      RECT 1169.500000 294.350000 1170.500000 295.650000 ;
      RECT 1116.500000 294.350000 1149.500000 295.650000 ;
      RECT 1107.500000 294.350000 1108.500000 295.650000 ;
      RECT 1066.500000 294.350000 1099.500000 295.650000 ;
      RECT 1057.500000 294.350000 1058.500000 295.650000 ;
      RECT 1016.500000 294.350000 1049.500000 295.650000 ;
      RECT 1007.500000 294.350000 1008.500000 295.650000 ;
      RECT 966.500000 294.350000 999.500000 295.650000 ;
      RECT 957.500000 294.350000 958.500000 295.650000 ;
      RECT 916.500000 294.350000 949.500000 295.650000 ;
      RECT 907.500000 294.350000 908.500000 295.650000 ;
      RECT 866.500000 294.350000 899.500000 295.650000 ;
      RECT 857.500000 294.350000 858.500000 295.650000 ;
      RECT 816.500000 294.350000 849.500000 295.650000 ;
      RECT 807.500000 294.350000 808.500000 295.650000 ;
      RECT 766.500000 294.350000 799.500000 295.650000 ;
      RECT 757.500000 294.350000 758.500000 295.650000 ;
      RECT 716.500000 294.350000 749.500000 295.650000 ;
      RECT 707.500000 294.350000 708.500000 295.650000 ;
      RECT 666.500000 294.350000 699.500000 295.650000 ;
      RECT 657.500000 294.350000 658.500000 295.650000 ;
      RECT 616.500000 294.350000 649.500000 295.650000 ;
      RECT 607.500000 294.350000 608.500000 295.650000 ;
      RECT 566.500000 294.350000 599.500000 295.650000 ;
      RECT 557.500000 294.350000 558.500000 295.650000 ;
      RECT 516.500000 294.350000 549.500000 295.650000 ;
      RECT 507.500000 294.350000 508.500000 295.650000 ;
      RECT 466.500000 294.350000 499.500000 295.650000 ;
      RECT 457.500000 294.350000 458.500000 295.650000 ;
      RECT 416.500000 294.350000 449.500000 295.650000 ;
      RECT 407.500000 294.350000 408.500000 295.650000 ;
      RECT 366.500000 294.350000 399.500000 295.650000 ;
      RECT 357.500000 294.350000 358.500000 295.650000 ;
      RECT 316.500000 294.350000 349.500000 295.650000 ;
      RECT 307.500000 294.350000 308.500000 295.650000 ;
      RECT 266.500000 294.350000 299.500000 295.650000 ;
      RECT 257.500000 294.350000 258.500000 295.650000 ;
      RECT 216.500000 294.350000 249.500000 295.650000 ;
      RECT 207.500000 294.350000 208.500000 295.650000 ;
      RECT 166.500000 294.350000 199.500000 295.650000 ;
      RECT 157.500000 294.350000 158.500000 295.650000 ;
      RECT 116.500000 294.350000 149.500000 295.650000 ;
      RECT 107.500000 294.350000 108.500000 295.650000 ;
      RECT 66.500000 294.350000 99.500000 295.650000 ;
      RECT 57.500000 294.350000 58.500000 295.650000 ;
      RECT 29.500000 294.350000 49.500000 295.650000 ;
      RECT 15.500000 294.350000 16.500000 295.650000 ;
      RECT 1157.500000 293.650000 1170.500000 294.350000 ;
      RECT 1107.500000 293.650000 1149.500000 294.350000 ;
      RECT 1057.500000 293.650000 1099.500000 294.350000 ;
      RECT 1007.500000 293.650000 1049.500000 294.350000 ;
      RECT 957.500000 293.650000 999.500000 294.350000 ;
      RECT 907.500000 293.650000 949.500000 294.350000 ;
      RECT 857.500000 293.650000 899.500000 294.350000 ;
      RECT 807.500000 293.650000 849.500000 294.350000 ;
      RECT 757.500000 293.650000 799.500000 294.350000 ;
      RECT 707.500000 293.650000 749.500000 294.350000 ;
      RECT 657.500000 293.650000 699.500000 294.350000 ;
      RECT 607.500000 293.650000 649.500000 294.350000 ;
      RECT 557.500000 293.650000 599.500000 294.350000 ;
      RECT 507.500000 293.650000 549.500000 294.350000 ;
      RECT 457.500000 293.650000 499.500000 294.350000 ;
      RECT 407.500000 293.650000 449.500000 294.350000 ;
      RECT 357.500000 293.650000 399.500000 294.350000 ;
      RECT 307.500000 293.650000 349.500000 294.350000 ;
      RECT 257.500000 293.650000 299.500000 294.350000 ;
      RECT 207.500000 293.650000 249.500000 294.350000 ;
      RECT 157.500000 293.650000 199.500000 294.350000 ;
      RECT 107.500000 293.650000 149.500000 294.350000 ;
      RECT 57.500000 293.650000 99.500000 294.350000 ;
      RECT 15.500000 293.650000 49.500000 294.350000 ;
      RECT 2.020000 293.515000 2.500000 295.650000 ;
      RECT 1183.500000 292.350000 1186.000000 295.650000 ;
      RECT 1169.500000 292.350000 1170.500000 293.650000 ;
      RECT 1116.500000 292.350000 1149.500000 293.650000 ;
      RECT 1107.500000 292.350000 1108.500000 293.650000 ;
      RECT 1066.500000 292.350000 1099.500000 293.650000 ;
      RECT 1057.500000 292.350000 1058.500000 293.650000 ;
      RECT 1016.500000 292.350000 1049.500000 293.650000 ;
      RECT 1007.500000 292.350000 1008.500000 293.650000 ;
      RECT 966.500000 292.350000 999.500000 293.650000 ;
      RECT 957.500000 292.350000 958.500000 293.650000 ;
      RECT 916.500000 292.350000 949.500000 293.650000 ;
      RECT 907.500000 292.350000 908.500000 293.650000 ;
      RECT 866.500000 292.350000 899.500000 293.650000 ;
      RECT 857.500000 292.350000 858.500000 293.650000 ;
      RECT 816.500000 292.350000 849.500000 293.650000 ;
      RECT 807.500000 292.350000 808.500000 293.650000 ;
      RECT 766.500000 292.350000 799.500000 293.650000 ;
      RECT 757.500000 292.350000 758.500000 293.650000 ;
      RECT 716.500000 292.350000 749.500000 293.650000 ;
      RECT 707.500000 292.350000 708.500000 293.650000 ;
      RECT 666.500000 292.350000 699.500000 293.650000 ;
      RECT 657.500000 292.350000 658.500000 293.650000 ;
      RECT 616.500000 292.350000 649.500000 293.650000 ;
      RECT 607.500000 292.350000 608.500000 293.650000 ;
      RECT 566.500000 292.350000 599.500000 293.650000 ;
      RECT 557.500000 292.350000 558.500000 293.650000 ;
      RECT 516.500000 292.350000 549.500000 293.650000 ;
      RECT 507.500000 292.350000 508.500000 293.650000 ;
      RECT 466.500000 292.350000 499.500000 293.650000 ;
      RECT 457.500000 292.350000 458.500000 293.650000 ;
      RECT 416.500000 292.350000 449.500000 293.650000 ;
      RECT 407.500000 292.350000 408.500000 293.650000 ;
      RECT 366.500000 292.350000 399.500000 293.650000 ;
      RECT 357.500000 292.350000 358.500000 293.650000 ;
      RECT 316.500000 292.350000 349.500000 293.650000 ;
      RECT 307.500000 292.350000 308.500000 293.650000 ;
      RECT 266.500000 292.350000 299.500000 293.650000 ;
      RECT 257.500000 292.350000 258.500000 293.650000 ;
      RECT 216.500000 292.350000 249.500000 293.650000 ;
      RECT 207.500000 292.350000 208.500000 293.650000 ;
      RECT 166.500000 292.350000 199.500000 293.650000 ;
      RECT 157.500000 292.350000 158.500000 293.650000 ;
      RECT 116.500000 292.350000 149.500000 293.650000 ;
      RECT 107.500000 292.350000 108.500000 293.650000 ;
      RECT 66.500000 292.350000 99.500000 293.650000 ;
      RECT 57.500000 292.350000 58.500000 293.650000 ;
      RECT 29.500000 292.350000 49.500000 293.650000 ;
      RECT 15.500000 292.350000 16.500000 293.650000 ;
      RECT 0.000000 292.350000 2.500000 293.515000 ;
      RECT 1169.500000 291.650000 1186.000000 292.350000 ;
      RECT 1116.500000 291.650000 1156.500000 292.350000 ;
      RECT 1066.500000 291.650000 1108.500000 292.350000 ;
      RECT 1016.500000 291.650000 1058.500000 292.350000 ;
      RECT 966.500000 291.650000 1008.500000 292.350000 ;
      RECT 916.500000 291.650000 958.500000 292.350000 ;
      RECT 866.500000 291.650000 908.500000 292.350000 ;
      RECT 816.500000 291.650000 858.500000 292.350000 ;
      RECT 766.500000 291.650000 808.500000 292.350000 ;
      RECT 716.500000 291.650000 758.500000 292.350000 ;
      RECT 666.500000 291.650000 708.500000 292.350000 ;
      RECT 616.500000 291.650000 658.500000 292.350000 ;
      RECT 566.500000 291.650000 608.500000 292.350000 ;
      RECT 516.500000 291.650000 558.500000 292.350000 ;
      RECT 466.500000 291.650000 508.500000 292.350000 ;
      RECT 416.500000 291.650000 458.500000 292.350000 ;
      RECT 366.500000 291.650000 408.500000 292.350000 ;
      RECT 316.500000 291.650000 358.500000 292.350000 ;
      RECT 266.500000 291.650000 308.500000 292.350000 ;
      RECT 216.500000 291.650000 258.500000 292.350000 ;
      RECT 166.500000 291.650000 208.500000 292.350000 ;
      RECT 116.500000 291.650000 158.500000 292.350000 ;
      RECT 66.500000 291.650000 108.500000 292.350000 ;
      RECT 29.500000 291.650000 58.500000 292.350000 ;
      RECT 0.000000 291.650000 16.500000 292.350000 ;
      RECT 0.000000 290.935000 2.500000 291.650000 ;
      RECT 1183.500000 290.930000 1186.000000 291.650000 ;
      RECT 1169.500000 290.350000 1170.500000 291.650000 ;
      RECT 1116.500000 290.350000 1149.500000 291.650000 ;
      RECT 1107.500000 290.350000 1108.500000 291.650000 ;
      RECT 1066.500000 290.350000 1099.500000 291.650000 ;
      RECT 1057.500000 290.350000 1058.500000 291.650000 ;
      RECT 1016.500000 290.350000 1049.500000 291.650000 ;
      RECT 1007.500000 290.350000 1008.500000 291.650000 ;
      RECT 966.500000 290.350000 999.500000 291.650000 ;
      RECT 957.500000 290.350000 958.500000 291.650000 ;
      RECT 916.500000 290.350000 949.500000 291.650000 ;
      RECT 907.500000 290.350000 908.500000 291.650000 ;
      RECT 866.500000 290.350000 899.500000 291.650000 ;
      RECT 857.500000 290.350000 858.500000 291.650000 ;
      RECT 816.500000 290.350000 849.500000 291.650000 ;
      RECT 807.500000 290.350000 808.500000 291.650000 ;
      RECT 766.500000 290.350000 799.500000 291.650000 ;
      RECT 757.500000 290.350000 758.500000 291.650000 ;
      RECT 716.500000 290.350000 749.500000 291.650000 ;
      RECT 707.500000 290.350000 708.500000 291.650000 ;
      RECT 666.500000 290.350000 699.500000 291.650000 ;
      RECT 657.500000 290.350000 658.500000 291.650000 ;
      RECT 616.500000 290.350000 649.500000 291.650000 ;
      RECT 607.500000 290.350000 608.500000 291.650000 ;
      RECT 566.500000 290.350000 599.500000 291.650000 ;
      RECT 557.500000 290.350000 558.500000 291.650000 ;
      RECT 516.500000 290.350000 549.500000 291.650000 ;
      RECT 507.500000 290.350000 508.500000 291.650000 ;
      RECT 466.500000 290.350000 499.500000 291.650000 ;
      RECT 457.500000 290.350000 458.500000 291.650000 ;
      RECT 416.500000 290.350000 449.500000 291.650000 ;
      RECT 407.500000 290.350000 408.500000 291.650000 ;
      RECT 366.500000 290.350000 399.500000 291.650000 ;
      RECT 357.500000 290.350000 358.500000 291.650000 ;
      RECT 316.500000 290.350000 349.500000 291.650000 ;
      RECT 307.500000 290.350000 308.500000 291.650000 ;
      RECT 266.500000 290.350000 299.500000 291.650000 ;
      RECT 257.500000 290.350000 258.500000 291.650000 ;
      RECT 216.500000 290.350000 249.500000 291.650000 ;
      RECT 207.500000 290.350000 208.500000 291.650000 ;
      RECT 166.500000 290.350000 199.500000 291.650000 ;
      RECT 157.500000 290.350000 158.500000 291.650000 ;
      RECT 116.500000 290.350000 149.500000 291.650000 ;
      RECT 107.500000 290.350000 108.500000 291.650000 ;
      RECT 66.500000 290.350000 99.500000 291.650000 ;
      RECT 57.500000 290.350000 58.500000 291.650000 ;
      RECT 29.500000 290.350000 49.500000 291.650000 ;
      RECT 15.500000 290.350000 16.500000 291.650000 ;
      RECT 1157.500000 289.650000 1170.500000 290.350000 ;
      RECT 1107.500000 289.650000 1149.500000 290.350000 ;
      RECT 1057.500000 289.650000 1099.500000 290.350000 ;
      RECT 1007.500000 289.650000 1049.500000 290.350000 ;
      RECT 957.500000 289.650000 999.500000 290.350000 ;
      RECT 907.500000 289.650000 949.500000 290.350000 ;
      RECT 857.500000 289.650000 899.500000 290.350000 ;
      RECT 807.500000 289.650000 849.500000 290.350000 ;
      RECT 757.500000 289.650000 799.500000 290.350000 ;
      RECT 707.500000 289.650000 749.500000 290.350000 ;
      RECT 657.500000 289.650000 699.500000 290.350000 ;
      RECT 607.500000 289.650000 649.500000 290.350000 ;
      RECT 557.500000 289.650000 599.500000 290.350000 ;
      RECT 507.500000 289.650000 549.500000 290.350000 ;
      RECT 457.500000 289.650000 499.500000 290.350000 ;
      RECT 407.500000 289.650000 449.500000 290.350000 ;
      RECT 357.500000 289.650000 399.500000 290.350000 ;
      RECT 307.500000 289.650000 349.500000 290.350000 ;
      RECT 257.500000 289.650000 299.500000 290.350000 ;
      RECT 207.500000 289.650000 249.500000 290.350000 ;
      RECT 157.500000 289.650000 199.500000 290.350000 ;
      RECT 107.500000 289.650000 149.500000 290.350000 ;
      RECT 57.500000 289.650000 99.500000 290.350000 ;
      RECT 15.500000 289.650000 49.500000 290.350000 ;
      RECT 1183.500000 288.350000 1183.980000 290.930000 ;
      RECT 1169.500000 288.350000 1170.500000 289.650000 ;
      RECT 1116.500000 288.350000 1149.500000 289.650000 ;
      RECT 1107.500000 288.350000 1108.500000 289.650000 ;
      RECT 1066.500000 288.350000 1099.500000 289.650000 ;
      RECT 1057.500000 288.350000 1058.500000 289.650000 ;
      RECT 1016.500000 288.350000 1049.500000 289.650000 ;
      RECT 1007.500000 288.350000 1008.500000 289.650000 ;
      RECT 966.500000 288.350000 999.500000 289.650000 ;
      RECT 957.500000 288.350000 958.500000 289.650000 ;
      RECT 916.500000 288.350000 949.500000 289.650000 ;
      RECT 907.500000 288.350000 908.500000 289.650000 ;
      RECT 866.500000 288.350000 899.500000 289.650000 ;
      RECT 857.500000 288.350000 858.500000 289.650000 ;
      RECT 816.500000 288.350000 849.500000 289.650000 ;
      RECT 807.500000 288.350000 808.500000 289.650000 ;
      RECT 766.500000 288.350000 799.500000 289.650000 ;
      RECT 757.500000 288.350000 758.500000 289.650000 ;
      RECT 716.500000 288.350000 749.500000 289.650000 ;
      RECT 707.500000 288.350000 708.500000 289.650000 ;
      RECT 666.500000 288.350000 699.500000 289.650000 ;
      RECT 657.500000 288.350000 658.500000 289.650000 ;
      RECT 616.500000 288.350000 649.500000 289.650000 ;
      RECT 607.500000 288.350000 608.500000 289.650000 ;
      RECT 566.500000 288.350000 599.500000 289.650000 ;
      RECT 557.500000 288.350000 558.500000 289.650000 ;
      RECT 516.500000 288.350000 549.500000 289.650000 ;
      RECT 507.500000 288.350000 508.500000 289.650000 ;
      RECT 466.500000 288.350000 499.500000 289.650000 ;
      RECT 457.500000 288.350000 458.500000 289.650000 ;
      RECT 416.500000 288.350000 449.500000 289.650000 ;
      RECT 407.500000 288.350000 408.500000 289.650000 ;
      RECT 366.500000 288.350000 399.500000 289.650000 ;
      RECT 357.500000 288.350000 358.500000 289.650000 ;
      RECT 316.500000 288.350000 349.500000 289.650000 ;
      RECT 307.500000 288.350000 308.500000 289.650000 ;
      RECT 266.500000 288.350000 299.500000 289.650000 ;
      RECT 257.500000 288.350000 258.500000 289.650000 ;
      RECT 216.500000 288.350000 249.500000 289.650000 ;
      RECT 207.500000 288.350000 208.500000 289.650000 ;
      RECT 166.500000 288.350000 199.500000 289.650000 ;
      RECT 157.500000 288.350000 158.500000 289.650000 ;
      RECT 116.500000 288.350000 149.500000 289.650000 ;
      RECT 107.500000 288.350000 108.500000 289.650000 ;
      RECT 66.500000 288.350000 99.500000 289.650000 ;
      RECT 57.500000 288.350000 58.500000 289.650000 ;
      RECT 29.500000 288.350000 49.500000 289.650000 ;
      RECT 15.500000 288.350000 16.500000 289.650000 ;
      RECT 2.020000 288.350000 2.500000 290.935000 ;
      RECT 2.020000 287.835000 16.500000 288.350000 ;
      RECT 1169.500000 287.830000 1183.980000 288.350000 ;
      RECT 1169.500000 287.650000 1186.000000 287.830000 ;
      RECT 1116.500000 287.650000 1156.500000 288.350000 ;
      RECT 1066.500000 287.650000 1108.500000 288.350000 ;
      RECT 1016.500000 287.650000 1058.500000 288.350000 ;
      RECT 966.500000 287.650000 1008.500000 288.350000 ;
      RECT 916.500000 287.650000 958.500000 288.350000 ;
      RECT 866.500000 287.650000 908.500000 288.350000 ;
      RECT 816.500000 287.650000 858.500000 288.350000 ;
      RECT 766.500000 287.650000 808.500000 288.350000 ;
      RECT 716.500000 287.650000 758.500000 288.350000 ;
      RECT 666.500000 287.650000 708.500000 288.350000 ;
      RECT 616.500000 287.650000 658.500000 288.350000 ;
      RECT 566.500000 287.650000 608.500000 288.350000 ;
      RECT 516.500000 287.650000 558.500000 288.350000 ;
      RECT 466.500000 287.650000 508.500000 288.350000 ;
      RECT 416.500000 287.650000 458.500000 288.350000 ;
      RECT 366.500000 287.650000 408.500000 288.350000 ;
      RECT 316.500000 287.650000 358.500000 288.350000 ;
      RECT 266.500000 287.650000 308.500000 288.350000 ;
      RECT 216.500000 287.650000 258.500000 288.350000 ;
      RECT 166.500000 287.650000 208.500000 288.350000 ;
      RECT 116.500000 287.650000 158.500000 288.350000 ;
      RECT 66.500000 287.650000 108.500000 288.350000 ;
      RECT 29.500000 287.650000 58.500000 288.350000 ;
      RECT 0.000000 287.650000 16.500000 287.835000 ;
      RECT 1169.500000 286.350000 1170.500000 287.650000 ;
      RECT 1116.500000 286.350000 1149.500000 287.650000 ;
      RECT 1107.500000 286.350000 1108.500000 287.650000 ;
      RECT 1066.500000 286.350000 1099.500000 287.650000 ;
      RECT 1057.500000 286.350000 1058.500000 287.650000 ;
      RECT 1016.500000 286.350000 1049.500000 287.650000 ;
      RECT 1007.500000 286.350000 1008.500000 287.650000 ;
      RECT 966.500000 286.350000 999.500000 287.650000 ;
      RECT 957.500000 286.350000 958.500000 287.650000 ;
      RECT 916.500000 286.350000 949.500000 287.650000 ;
      RECT 907.500000 286.350000 908.500000 287.650000 ;
      RECT 866.500000 286.350000 899.500000 287.650000 ;
      RECT 857.500000 286.350000 858.500000 287.650000 ;
      RECT 816.500000 286.350000 849.500000 287.650000 ;
      RECT 807.500000 286.350000 808.500000 287.650000 ;
      RECT 766.500000 286.350000 799.500000 287.650000 ;
      RECT 757.500000 286.350000 758.500000 287.650000 ;
      RECT 716.500000 286.350000 749.500000 287.650000 ;
      RECT 707.500000 286.350000 708.500000 287.650000 ;
      RECT 666.500000 286.350000 699.500000 287.650000 ;
      RECT 657.500000 286.350000 658.500000 287.650000 ;
      RECT 616.500000 286.350000 649.500000 287.650000 ;
      RECT 607.500000 286.350000 608.500000 287.650000 ;
      RECT 566.500000 286.350000 599.500000 287.650000 ;
      RECT 557.500000 286.350000 558.500000 287.650000 ;
      RECT 516.500000 286.350000 549.500000 287.650000 ;
      RECT 507.500000 286.350000 508.500000 287.650000 ;
      RECT 466.500000 286.350000 499.500000 287.650000 ;
      RECT 457.500000 286.350000 458.500000 287.650000 ;
      RECT 416.500000 286.350000 449.500000 287.650000 ;
      RECT 407.500000 286.350000 408.500000 287.650000 ;
      RECT 366.500000 286.350000 399.500000 287.650000 ;
      RECT 357.500000 286.350000 358.500000 287.650000 ;
      RECT 316.500000 286.350000 349.500000 287.650000 ;
      RECT 307.500000 286.350000 308.500000 287.650000 ;
      RECT 266.500000 286.350000 299.500000 287.650000 ;
      RECT 257.500000 286.350000 258.500000 287.650000 ;
      RECT 216.500000 286.350000 249.500000 287.650000 ;
      RECT 207.500000 286.350000 208.500000 287.650000 ;
      RECT 166.500000 286.350000 199.500000 287.650000 ;
      RECT 157.500000 286.350000 158.500000 287.650000 ;
      RECT 116.500000 286.350000 149.500000 287.650000 ;
      RECT 107.500000 286.350000 108.500000 287.650000 ;
      RECT 66.500000 286.350000 99.500000 287.650000 ;
      RECT 57.500000 286.350000 58.500000 287.650000 ;
      RECT 29.500000 286.350000 49.500000 287.650000 ;
      RECT 15.500000 286.350000 16.500000 287.650000 ;
      RECT 1157.500000 285.650000 1170.500000 286.350000 ;
      RECT 1107.500000 285.650000 1149.500000 286.350000 ;
      RECT 1057.500000 285.650000 1099.500000 286.350000 ;
      RECT 1007.500000 285.650000 1049.500000 286.350000 ;
      RECT 957.500000 285.650000 999.500000 286.350000 ;
      RECT 907.500000 285.650000 949.500000 286.350000 ;
      RECT 857.500000 285.650000 899.500000 286.350000 ;
      RECT 807.500000 285.650000 849.500000 286.350000 ;
      RECT 757.500000 285.650000 799.500000 286.350000 ;
      RECT 707.500000 285.650000 749.500000 286.350000 ;
      RECT 657.500000 285.650000 699.500000 286.350000 ;
      RECT 607.500000 285.650000 649.500000 286.350000 ;
      RECT 557.500000 285.650000 599.500000 286.350000 ;
      RECT 507.500000 285.650000 549.500000 286.350000 ;
      RECT 457.500000 285.650000 499.500000 286.350000 ;
      RECT 407.500000 285.650000 449.500000 286.350000 ;
      RECT 357.500000 285.650000 399.500000 286.350000 ;
      RECT 307.500000 285.650000 349.500000 286.350000 ;
      RECT 257.500000 285.650000 299.500000 286.350000 ;
      RECT 207.500000 285.650000 249.500000 286.350000 ;
      RECT 157.500000 285.650000 199.500000 286.350000 ;
      RECT 107.500000 285.650000 149.500000 286.350000 ;
      RECT 57.500000 285.650000 99.500000 286.350000 ;
      RECT 15.500000 285.650000 49.500000 286.350000 ;
      RECT 1183.500000 284.350000 1186.000000 287.650000 ;
      RECT 1169.500000 284.350000 1170.500000 285.650000 ;
      RECT 1116.500000 284.350000 1149.500000 285.650000 ;
      RECT 1107.500000 284.350000 1108.500000 285.650000 ;
      RECT 1066.500000 284.350000 1099.500000 285.650000 ;
      RECT 1057.500000 284.350000 1058.500000 285.650000 ;
      RECT 1016.500000 284.350000 1049.500000 285.650000 ;
      RECT 1007.500000 284.350000 1008.500000 285.650000 ;
      RECT 966.500000 284.350000 999.500000 285.650000 ;
      RECT 957.500000 284.350000 958.500000 285.650000 ;
      RECT 916.500000 284.350000 949.500000 285.650000 ;
      RECT 907.500000 284.350000 908.500000 285.650000 ;
      RECT 866.500000 284.350000 899.500000 285.650000 ;
      RECT 857.500000 284.350000 858.500000 285.650000 ;
      RECT 816.500000 284.350000 849.500000 285.650000 ;
      RECT 807.500000 284.350000 808.500000 285.650000 ;
      RECT 766.500000 284.350000 799.500000 285.650000 ;
      RECT 757.500000 284.350000 758.500000 285.650000 ;
      RECT 716.500000 284.350000 749.500000 285.650000 ;
      RECT 707.500000 284.350000 708.500000 285.650000 ;
      RECT 666.500000 284.350000 699.500000 285.650000 ;
      RECT 657.500000 284.350000 658.500000 285.650000 ;
      RECT 616.500000 284.350000 649.500000 285.650000 ;
      RECT 607.500000 284.350000 608.500000 285.650000 ;
      RECT 566.500000 284.350000 599.500000 285.650000 ;
      RECT 557.500000 284.350000 558.500000 285.650000 ;
      RECT 516.500000 284.350000 549.500000 285.650000 ;
      RECT 507.500000 284.350000 508.500000 285.650000 ;
      RECT 466.500000 284.350000 499.500000 285.650000 ;
      RECT 457.500000 284.350000 458.500000 285.650000 ;
      RECT 416.500000 284.350000 449.500000 285.650000 ;
      RECT 407.500000 284.350000 408.500000 285.650000 ;
      RECT 366.500000 284.350000 399.500000 285.650000 ;
      RECT 357.500000 284.350000 358.500000 285.650000 ;
      RECT 316.500000 284.350000 349.500000 285.650000 ;
      RECT 307.500000 284.350000 308.500000 285.650000 ;
      RECT 266.500000 284.350000 299.500000 285.650000 ;
      RECT 257.500000 284.350000 258.500000 285.650000 ;
      RECT 216.500000 284.350000 249.500000 285.650000 ;
      RECT 207.500000 284.350000 208.500000 285.650000 ;
      RECT 166.500000 284.350000 199.500000 285.650000 ;
      RECT 157.500000 284.350000 158.500000 285.650000 ;
      RECT 116.500000 284.350000 149.500000 285.650000 ;
      RECT 107.500000 284.350000 108.500000 285.650000 ;
      RECT 66.500000 284.350000 99.500000 285.650000 ;
      RECT 57.500000 284.350000 58.500000 285.650000 ;
      RECT 29.500000 284.350000 49.500000 285.650000 ;
      RECT 15.500000 284.350000 16.500000 285.650000 ;
      RECT 0.000000 284.350000 2.500000 287.650000 ;
      RECT 1169.500000 283.650000 1186.000000 284.350000 ;
      RECT 1116.500000 283.650000 1156.500000 284.350000 ;
      RECT 1066.500000 283.650000 1108.500000 284.350000 ;
      RECT 1016.500000 283.650000 1058.500000 284.350000 ;
      RECT 966.500000 283.650000 1008.500000 284.350000 ;
      RECT 916.500000 283.650000 958.500000 284.350000 ;
      RECT 866.500000 283.650000 908.500000 284.350000 ;
      RECT 816.500000 283.650000 858.500000 284.350000 ;
      RECT 766.500000 283.650000 808.500000 284.350000 ;
      RECT 716.500000 283.650000 758.500000 284.350000 ;
      RECT 666.500000 283.650000 708.500000 284.350000 ;
      RECT 616.500000 283.650000 658.500000 284.350000 ;
      RECT 566.500000 283.650000 608.500000 284.350000 ;
      RECT 516.500000 283.650000 558.500000 284.350000 ;
      RECT 466.500000 283.650000 508.500000 284.350000 ;
      RECT 416.500000 283.650000 458.500000 284.350000 ;
      RECT 366.500000 283.650000 408.500000 284.350000 ;
      RECT 316.500000 283.650000 358.500000 284.350000 ;
      RECT 266.500000 283.650000 308.500000 284.350000 ;
      RECT 216.500000 283.650000 258.500000 284.350000 ;
      RECT 166.500000 283.650000 208.500000 284.350000 ;
      RECT 116.500000 283.650000 158.500000 284.350000 ;
      RECT 66.500000 283.650000 108.500000 284.350000 ;
      RECT 29.500000 283.650000 58.500000 284.350000 ;
      RECT 0.000000 283.650000 16.500000 284.350000 ;
      RECT 1169.500000 282.350000 1170.500000 283.650000 ;
      RECT 1116.500000 282.350000 1149.500000 283.650000 ;
      RECT 1107.500000 282.350000 1108.500000 283.650000 ;
      RECT 1066.500000 282.350000 1099.500000 283.650000 ;
      RECT 1057.500000 282.350000 1058.500000 283.650000 ;
      RECT 1016.500000 282.350000 1049.500000 283.650000 ;
      RECT 1007.500000 282.350000 1008.500000 283.650000 ;
      RECT 966.500000 282.350000 999.500000 283.650000 ;
      RECT 957.500000 282.350000 958.500000 283.650000 ;
      RECT 916.500000 282.350000 949.500000 283.650000 ;
      RECT 907.500000 282.350000 908.500000 283.650000 ;
      RECT 866.500000 282.350000 899.500000 283.650000 ;
      RECT 857.500000 282.350000 858.500000 283.650000 ;
      RECT 816.500000 282.350000 849.500000 283.650000 ;
      RECT 807.500000 282.350000 808.500000 283.650000 ;
      RECT 766.500000 282.350000 799.500000 283.650000 ;
      RECT 757.500000 282.350000 758.500000 283.650000 ;
      RECT 716.500000 282.350000 749.500000 283.650000 ;
      RECT 707.500000 282.350000 708.500000 283.650000 ;
      RECT 666.500000 282.350000 699.500000 283.650000 ;
      RECT 657.500000 282.350000 658.500000 283.650000 ;
      RECT 616.500000 282.350000 649.500000 283.650000 ;
      RECT 607.500000 282.350000 608.500000 283.650000 ;
      RECT 566.500000 282.350000 599.500000 283.650000 ;
      RECT 557.500000 282.350000 558.500000 283.650000 ;
      RECT 516.500000 282.350000 549.500000 283.650000 ;
      RECT 507.500000 282.350000 508.500000 283.650000 ;
      RECT 466.500000 282.350000 499.500000 283.650000 ;
      RECT 457.500000 282.350000 458.500000 283.650000 ;
      RECT 416.500000 282.350000 449.500000 283.650000 ;
      RECT 407.500000 282.350000 408.500000 283.650000 ;
      RECT 366.500000 282.350000 399.500000 283.650000 ;
      RECT 357.500000 282.350000 358.500000 283.650000 ;
      RECT 316.500000 282.350000 349.500000 283.650000 ;
      RECT 307.500000 282.350000 308.500000 283.650000 ;
      RECT 266.500000 282.350000 299.500000 283.650000 ;
      RECT 257.500000 282.350000 258.500000 283.650000 ;
      RECT 216.500000 282.350000 249.500000 283.650000 ;
      RECT 207.500000 282.350000 208.500000 283.650000 ;
      RECT 166.500000 282.350000 199.500000 283.650000 ;
      RECT 157.500000 282.350000 158.500000 283.650000 ;
      RECT 116.500000 282.350000 149.500000 283.650000 ;
      RECT 107.500000 282.350000 108.500000 283.650000 ;
      RECT 66.500000 282.350000 99.500000 283.650000 ;
      RECT 57.500000 282.350000 58.500000 283.650000 ;
      RECT 29.500000 282.350000 49.500000 283.650000 ;
      RECT 15.500000 282.350000 16.500000 283.650000 ;
      RECT 1157.500000 281.650000 1170.500000 282.350000 ;
      RECT 1107.500000 281.650000 1149.500000 282.350000 ;
      RECT 1057.500000 281.650000 1099.500000 282.350000 ;
      RECT 1007.500000 281.650000 1049.500000 282.350000 ;
      RECT 957.500000 281.650000 999.500000 282.350000 ;
      RECT 907.500000 281.650000 949.500000 282.350000 ;
      RECT 857.500000 281.650000 899.500000 282.350000 ;
      RECT 807.500000 281.650000 849.500000 282.350000 ;
      RECT 757.500000 281.650000 799.500000 282.350000 ;
      RECT 707.500000 281.650000 749.500000 282.350000 ;
      RECT 657.500000 281.650000 699.500000 282.350000 ;
      RECT 607.500000 281.650000 649.500000 282.350000 ;
      RECT 557.500000 281.650000 599.500000 282.350000 ;
      RECT 507.500000 281.650000 549.500000 282.350000 ;
      RECT 457.500000 281.650000 499.500000 282.350000 ;
      RECT 407.500000 281.650000 449.500000 282.350000 ;
      RECT 357.500000 281.650000 399.500000 282.350000 ;
      RECT 307.500000 281.650000 349.500000 282.350000 ;
      RECT 257.500000 281.650000 299.500000 282.350000 ;
      RECT 207.500000 281.650000 249.500000 282.350000 ;
      RECT 157.500000 281.650000 199.500000 282.350000 ;
      RECT 107.500000 281.650000 149.500000 282.350000 ;
      RECT 57.500000 281.650000 99.500000 282.350000 ;
      RECT 15.500000 281.650000 49.500000 282.350000 ;
      RECT 1183.500000 280.350000 1186.000000 283.650000 ;
      RECT 1169.500000 280.350000 1170.500000 281.650000 ;
      RECT 1116.500000 280.350000 1149.500000 281.650000 ;
      RECT 1107.500000 280.350000 1108.500000 281.650000 ;
      RECT 1066.500000 280.350000 1099.500000 281.650000 ;
      RECT 1057.500000 280.350000 1058.500000 281.650000 ;
      RECT 1016.500000 280.350000 1049.500000 281.650000 ;
      RECT 1007.500000 280.350000 1008.500000 281.650000 ;
      RECT 966.500000 280.350000 999.500000 281.650000 ;
      RECT 957.500000 280.350000 958.500000 281.650000 ;
      RECT 916.500000 280.350000 949.500000 281.650000 ;
      RECT 907.500000 280.350000 908.500000 281.650000 ;
      RECT 866.500000 280.350000 899.500000 281.650000 ;
      RECT 857.500000 280.350000 858.500000 281.650000 ;
      RECT 816.500000 280.350000 849.500000 281.650000 ;
      RECT 807.500000 280.350000 808.500000 281.650000 ;
      RECT 766.500000 280.350000 799.500000 281.650000 ;
      RECT 757.500000 280.350000 758.500000 281.650000 ;
      RECT 716.500000 280.350000 749.500000 281.650000 ;
      RECT 707.500000 280.350000 708.500000 281.650000 ;
      RECT 666.500000 280.350000 699.500000 281.650000 ;
      RECT 657.500000 280.350000 658.500000 281.650000 ;
      RECT 616.500000 280.350000 649.500000 281.650000 ;
      RECT 607.500000 280.350000 608.500000 281.650000 ;
      RECT 566.500000 280.350000 599.500000 281.650000 ;
      RECT 557.500000 280.350000 558.500000 281.650000 ;
      RECT 516.500000 280.350000 549.500000 281.650000 ;
      RECT 507.500000 280.350000 508.500000 281.650000 ;
      RECT 466.500000 280.350000 499.500000 281.650000 ;
      RECT 457.500000 280.350000 458.500000 281.650000 ;
      RECT 416.500000 280.350000 449.500000 281.650000 ;
      RECT 407.500000 280.350000 408.500000 281.650000 ;
      RECT 366.500000 280.350000 399.500000 281.650000 ;
      RECT 357.500000 280.350000 358.500000 281.650000 ;
      RECT 316.500000 280.350000 349.500000 281.650000 ;
      RECT 307.500000 280.350000 308.500000 281.650000 ;
      RECT 266.500000 280.350000 299.500000 281.650000 ;
      RECT 257.500000 280.350000 258.500000 281.650000 ;
      RECT 216.500000 280.350000 249.500000 281.650000 ;
      RECT 207.500000 280.350000 208.500000 281.650000 ;
      RECT 166.500000 280.350000 199.500000 281.650000 ;
      RECT 157.500000 280.350000 158.500000 281.650000 ;
      RECT 116.500000 280.350000 149.500000 281.650000 ;
      RECT 107.500000 280.350000 108.500000 281.650000 ;
      RECT 66.500000 280.350000 99.500000 281.650000 ;
      RECT 57.500000 280.350000 58.500000 281.650000 ;
      RECT 29.500000 280.350000 49.500000 281.650000 ;
      RECT 15.500000 280.350000 16.500000 281.650000 ;
      RECT 0.000000 280.350000 2.500000 283.650000 ;
      RECT 1169.500000 279.650000 1186.000000 280.350000 ;
      RECT 1116.500000 279.650000 1156.500000 280.350000 ;
      RECT 1066.500000 279.650000 1108.500000 280.350000 ;
      RECT 1016.500000 279.650000 1058.500000 280.350000 ;
      RECT 966.500000 279.650000 1008.500000 280.350000 ;
      RECT 916.500000 279.650000 958.500000 280.350000 ;
      RECT 866.500000 279.650000 908.500000 280.350000 ;
      RECT 816.500000 279.650000 858.500000 280.350000 ;
      RECT 766.500000 279.650000 808.500000 280.350000 ;
      RECT 716.500000 279.650000 758.500000 280.350000 ;
      RECT 666.500000 279.650000 708.500000 280.350000 ;
      RECT 616.500000 279.650000 658.500000 280.350000 ;
      RECT 566.500000 279.650000 608.500000 280.350000 ;
      RECT 516.500000 279.650000 558.500000 280.350000 ;
      RECT 466.500000 279.650000 508.500000 280.350000 ;
      RECT 416.500000 279.650000 458.500000 280.350000 ;
      RECT 366.500000 279.650000 408.500000 280.350000 ;
      RECT 316.500000 279.650000 358.500000 280.350000 ;
      RECT 266.500000 279.650000 308.500000 280.350000 ;
      RECT 216.500000 279.650000 258.500000 280.350000 ;
      RECT 166.500000 279.650000 208.500000 280.350000 ;
      RECT 116.500000 279.650000 158.500000 280.350000 ;
      RECT 66.500000 279.650000 108.500000 280.350000 ;
      RECT 29.500000 279.650000 58.500000 280.350000 ;
      RECT 0.000000 279.650000 16.500000 280.350000 ;
      RECT 1169.500000 278.350000 1170.500000 279.650000 ;
      RECT 1116.500000 278.350000 1149.500000 279.650000 ;
      RECT 1107.500000 278.350000 1108.500000 279.650000 ;
      RECT 1066.500000 278.350000 1099.500000 279.650000 ;
      RECT 1057.500000 278.350000 1058.500000 279.650000 ;
      RECT 1016.500000 278.350000 1049.500000 279.650000 ;
      RECT 1007.500000 278.350000 1008.500000 279.650000 ;
      RECT 966.500000 278.350000 999.500000 279.650000 ;
      RECT 957.500000 278.350000 958.500000 279.650000 ;
      RECT 916.500000 278.350000 949.500000 279.650000 ;
      RECT 907.500000 278.350000 908.500000 279.650000 ;
      RECT 866.500000 278.350000 899.500000 279.650000 ;
      RECT 857.500000 278.350000 858.500000 279.650000 ;
      RECT 816.500000 278.350000 849.500000 279.650000 ;
      RECT 807.500000 278.350000 808.500000 279.650000 ;
      RECT 766.500000 278.350000 799.500000 279.650000 ;
      RECT 757.500000 278.350000 758.500000 279.650000 ;
      RECT 716.500000 278.350000 749.500000 279.650000 ;
      RECT 707.500000 278.350000 708.500000 279.650000 ;
      RECT 666.500000 278.350000 699.500000 279.650000 ;
      RECT 657.500000 278.350000 658.500000 279.650000 ;
      RECT 616.500000 278.350000 649.500000 279.650000 ;
      RECT 607.500000 278.350000 608.500000 279.650000 ;
      RECT 566.500000 278.350000 599.500000 279.650000 ;
      RECT 557.500000 278.350000 558.500000 279.650000 ;
      RECT 516.500000 278.350000 549.500000 279.650000 ;
      RECT 507.500000 278.350000 508.500000 279.650000 ;
      RECT 466.500000 278.350000 499.500000 279.650000 ;
      RECT 457.500000 278.350000 458.500000 279.650000 ;
      RECT 416.500000 278.350000 449.500000 279.650000 ;
      RECT 407.500000 278.350000 408.500000 279.650000 ;
      RECT 366.500000 278.350000 399.500000 279.650000 ;
      RECT 357.500000 278.350000 358.500000 279.650000 ;
      RECT 316.500000 278.350000 349.500000 279.650000 ;
      RECT 307.500000 278.350000 308.500000 279.650000 ;
      RECT 266.500000 278.350000 299.500000 279.650000 ;
      RECT 257.500000 278.350000 258.500000 279.650000 ;
      RECT 216.500000 278.350000 249.500000 279.650000 ;
      RECT 207.500000 278.350000 208.500000 279.650000 ;
      RECT 166.500000 278.350000 199.500000 279.650000 ;
      RECT 157.500000 278.350000 158.500000 279.650000 ;
      RECT 116.500000 278.350000 149.500000 279.650000 ;
      RECT 107.500000 278.350000 108.500000 279.650000 ;
      RECT 66.500000 278.350000 99.500000 279.650000 ;
      RECT 57.500000 278.350000 58.500000 279.650000 ;
      RECT 29.500000 278.350000 49.500000 279.650000 ;
      RECT 15.500000 278.350000 16.500000 279.650000 ;
      RECT 1157.500000 277.650000 1170.500000 278.350000 ;
      RECT 1107.500000 277.650000 1149.500000 278.350000 ;
      RECT 1057.500000 277.650000 1099.500000 278.350000 ;
      RECT 1007.500000 277.650000 1049.500000 278.350000 ;
      RECT 957.500000 277.650000 999.500000 278.350000 ;
      RECT 907.500000 277.650000 949.500000 278.350000 ;
      RECT 857.500000 277.650000 899.500000 278.350000 ;
      RECT 807.500000 277.650000 849.500000 278.350000 ;
      RECT 757.500000 277.650000 799.500000 278.350000 ;
      RECT 707.500000 277.650000 749.500000 278.350000 ;
      RECT 657.500000 277.650000 699.500000 278.350000 ;
      RECT 607.500000 277.650000 649.500000 278.350000 ;
      RECT 557.500000 277.650000 599.500000 278.350000 ;
      RECT 507.500000 277.650000 549.500000 278.350000 ;
      RECT 457.500000 277.650000 499.500000 278.350000 ;
      RECT 407.500000 277.650000 449.500000 278.350000 ;
      RECT 357.500000 277.650000 399.500000 278.350000 ;
      RECT 307.500000 277.650000 349.500000 278.350000 ;
      RECT 257.500000 277.650000 299.500000 278.350000 ;
      RECT 207.500000 277.650000 249.500000 278.350000 ;
      RECT 157.500000 277.650000 199.500000 278.350000 ;
      RECT 107.500000 277.650000 149.500000 278.350000 ;
      RECT 57.500000 277.650000 99.500000 278.350000 ;
      RECT 15.500000 277.650000 49.500000 278.350000 ;
      RECT 1183.500000 276.350000 1186.000000 279.650000 ;
      RECT 1169.500000 276.350000 1170.500000 277.650000 ;
      RECT 1116.500000 276.350000 1149.500000 277.650000 ;
      RECT 1107.500000 276.350000 1108.500000 277.650000 ;
      RECT 1066.500000 276.350000 1099.500000 277.650000 ;
      RECT 1057.500000 276.350000 1058.500000 277.650000 ;
      RECT 1016.500000 276.350000 1049.500000 277.650000 ;
      RECT 1007.500000 276.350000 1008.500000 277.650000 ;
      RECT 966.500000 276.350000 999.500000 277.650000 ;
      RECT 957.500000 276.350000 958.500000 277.650000 ;
      RECT 916.500000 276.350000 949.500000 277.650000 ;
      RECT 907.500000 276.350000 908.500000 277.650000 ;
      RECT 866.500000 276.350000 899.500000 277.650000 ;
      RECT 857.500000 276.350000 858.500000 277.650000 ;
      RECT 816.500000 276.350000 849.500000 277.650000 ;
      RECT 807.500000 276.350000 808.500000 277.650000 ;
      RECT 766.500000 276.350000 799.500000 277.650000 ;
      RECT 757.500000 276.350000 758.500000 277.650000 ;
      RECT 716.500000 276.350000 749.500000 277.650000 ;
      RECT 707.500000 276.350000 708.500000 277.650000 ;
      RECT 666.500000 276.350000 699.500000 277.650000 ;
      RECT 657.500000 276.350000 658.500000 277.650000 ;
      RECT 616.500000 276.350000 649.500000 277.650000 ;
      RECT 607.500000 276.350000 608.500000 277.650000 ;
      RECT 566.500000 276.350000 599.500000 277.650000 ;
      RECT 557.500000 276.350000 558.500000 277.650000 ;
      RECT 516.500000 276.350000 549.500000 277.650000 ;
      RECT 507.500000 276.350000 508.500000 277.650000 ;
      RECT 466.500000 276.350000 499.500000 277.650000 ;
      RECT 457.500000 276.350000 458.500000 277.650000 ;
      RECT 416.500000 276.350000 449.500000 277.650000 ;
      RECT 407.500000 276.350000 408.500000 277.650000 ;
      RECT 366.500000 276.350000 399.500000 277.650000 ;
      RECT 357.500000 276.350000 358.500000 277.650000 ;
      RECT 316.500000 276.350000 349.500000 277.650000 ;
      RECT 307.500000 276.350000 308.500000 277.650000 ;
      RECT 266.500000 276.350000 299.500000 277.650000 ;
      RECT 257.500000 276.350000 258.500000 277.650000 ;
      RECT 216.500000 276.350000 249.500000 277.650000 ;
      RECT 207.500000 276.350000 208.500000 277.650000 ;
      RECT 166.500000 276.350000 199.500000 277.650000 ;
      RECT 157.500000 276.350000 158.500000 277.650000 ;
      RECT 116.500000 276.350000 149.500000 277.650000 ;
      RECT 107.500000 276.350000 108.500000 277.650000 ;
      RECT 66.500000 276.350000 99.500000 277.650000 ;
      RECT 57.500000 276.350000 58.500000 277.650000 ;
      RECT 29.500000 276.350000 49.500000 277.650000 ;
      RECT 15.500000 276.350000 16.500000 277.650000 ;
      RECT 0.000000 276.350000 2.500000 279.650000 ;
      RECT 1169.500000 275.650000 1186.000000 276.350000 ;
      RECT 1116.500000 275.650000 1156.500000 276.350000 ;
      RECT 1066.500000 275.650000 1108.500000 276.350000 ;
      RECT 1016.500000 275.650000 1058.500000 276.350000 ;
      RECT 966.500000 275.650000 1008.500000 276.350000 ;
      RECT 916.500000 275.650000 958.500000 276.350000 ;
      RECT 866.500000 275.650000 908.500000 276.350000 ;
      RECT 816.500000 275.650000 858.500000 276.350000 ;
      RECT 766.500000 275.650000 808.500000 276.350000 ;
      RECT 716.500000 275.650000 758.500000 276.350000 ;
      RECT 666.500000 275.650000 708.500000 276.350000 ;
      RECT 616.500000 275.650000 658.500000 276.350000 ;
      RECT 566.500000 275.650000 608.500000 276.350000 ;
      RECT 516.500000 275.650000 558.500000 276.350000 ;
      RECT 466.500000 275.650000 508.500000 276.350000 ;
      RECT 416.500000 275.650000 458.500000 276.350000 ;
      RECT 366.500000 275.650000 408.500000 276.350000 ;
      RECT 316.500000 275.650000 358.500000 276.350000 ;
      RECT 266.500000 275.650000 308.500000 276.350000 ;
      RECT 216.500000 275.650000 258.500000 276.350000 ;
      RECT 166.500000 275.650000 208.500000 276.350000 ;
      RECT 116.500000 275.650000 158.500000 276.350000 ;
      RECT 66.500000 275.650000 108.500000 276.350000 ;
      RECT 29.500000 275.650000 58.500000 276.350000 ;
      RECT 0.000000 275.650000 16.500000 276.350000 ;
      RECT 1169.500000 274.350000 1170.500000 275.650000 ;
      RECT 1116.500000 274.350000 1149.500000 275.650000 ;
      RECT 1107.500000 274.350000 1108.500000 275.650000 ;
      RECT 1066.500000 274.350000 1099.500000 275.650000 ;
      RECT 1057.500000 274.350000 1058.500000 275.650000 ;
      RECT 1016.500000 274.350000 1049.500000 275.650000 ;
      RECT 1007.500000 274.350000 1008.500000 275.650000 ;
      RECT 966.500000 274.350000 999.500000 275.650000 ;
      RECT 957.500000 274.350000 958.500000 275.650000 ;
      RECT 916.500000 274.350000 949.500000 275.650000 ;
      RECT 907.500000 274.350000 908.500000 275.650000 ;
      RECT 866.500000 274.350000 899.500000 275.650000 ;
      RECT 857.500000 274.350000 858.500000 275.650000 ;
      RECT 816.500000 274.350000 849.500000 275.650000 ;
      RECT 807.500000 274.350000 808.500000 275.650000 ;
      RECT 766.500000 274.350000 799.500000 275.650000 ;
      RECT 757.500000 274.350000 758.500000 275.650000 ;
      RECT 716.500000 274.350000 749.500000 275.650000 ;
      RECT 707.500000 274.350000 708.500000 275.650000 ;
      RECT 666.500000 274.350000 699.500000 275.650000 ;
      RECT 657.500000 274.350000 658.500000 275.650000 ;
      RECT 616.500000 274.350000 649.500000 275.650000 ;
      RECT 607.500000 274.350000 608.500000 275.650000 ;
      RECT 566.500000 274.350000 599.500000 275.650000 ;
      RECT 557.500000 274.350000 558.500000 275.650000 ;
      RECT 516.500000 274.350000 549.500000 275.650000 ;
      RECT 507.500000 274.350000 508.500000 275.650000 ;
      RECT 466.500000 274.350000 499.500000 275.650000 ;
      RECT 457.500000 274.350000 458.500000 275.650000 ;
      RECT 416.500000 274.350000 449.500000 275.650000 ;
      RECT 407.500000 274.350000 408.500000 275.650000 ;
      RECT 366.500000 274.350000 399.500000 275.650000 ;
      RECT 357.500000 274.350000 358.500000 275.650000 ;
      RECT 316.500000 274.350000 349.500000 275.650000 ;
      RECT 307.500000 274.350000 308.500000 275.650000 ;
      RECT 266.500000 274.350000 299.500000 275.650000 ;
      RECT 257.500000 274.350000 258.500000 275.650000 ;
      RECT 216.500000 274.350000 249.500000 275.650000 ;
      RECT 207.500000 274.350000 208.500000 275.650000 ;
      RECT 166.500000 274.350000 199.500000 275.650000 ;
      RECT 157.500000 274.350000 158.500000 275.650000 ;
      RECT 116.500000 274.350000 149.500000 275.650000 ;
      RECT 107.500000 274.350000 108.500000 275.650000 ;
      RECT 66.500000 274.350000 99.500000 275.650000 ;
      RECT 57.500000 274.350000 58.500000 275.650000 ;
      RECT 29.500000 274.350000 49.500000 275.650000 ;
      RECT 15.500000 274.350000 16.500000 275.650000 ;
      RECT 1157.500000 273.650000 1170.500000 274.350000 ;
      RECT 1107.500000 273.650000 1149.500000 274.350000 ;
      RECT 1057.500000 273.650000 1099.500000 274.350000 ;
      RECT 1007.500000 273.650000 1049.500000 274.350000 ;
      RECT 957.500000 273.650000 999.500000 274.350000 ;
      RECT 907.500000 273.650000 949.500000 274.350000 ;
      RECT 857.500000 273.650000 899.500000 274.350000 ;
      RECT 807.500000 273.650000 849.500000 274.350000 ;
      RECT 757.500000 273.650000 799.500000 274.350000 ;
      RECT 707.500000 273.650000 749.500000 274.350000 ;
      RECT 657.500000 273.650000 699.500000 274.350000 ;
      RECT 607.500000 273.650000 649.500000 274.350000 ;
      RECT 557.500000 273.650000 599.500000 274.350000 ;
      RECT 507.500000 273.650000 549.500000 274.350000 ;
      RECT 457.500000 273.650000 499.500000 274.350000 ;
      RECT 407.500000 273.650000 449.500000 274.350000 ;
      RECT 357.500000 273.650000 399.500000 274.350000 ;
      RECT 307.500000 273.650000 349.500000 274.350000 ;
      RECT 257.500000 273.650000 299.500000 274.350000 ;
      RECT 207.500000 273.650000 249.500000 274.350000 ;
      RECT 157.500000 273.650000 199.500000 274.350000 ;
      RECT 107.500000 273.650000 149.500000 274.350000 ;
      RECT 57.500000 273.650000 99.500000 274.350000 ;
      RECT 15.500000 273.650000 49.500000 274.350000 ;
      RECT 1183.500000 272.350000 1186.000000 275.650000 ;
      RECT 1169.500000 272.350000 1170.500000 273.650000 ;
      RECT 1116.500000 272.350000 1149.500000 273.650000 ;
      RECT 1107.500000 272.350000 1108.500000 273.650000 ;
      RECT 1066.500000 272.350000 1099.500000 273.650000 ;
      RECT 1057.500000 272.350000 1058.500000 273.650000 ;
      RECT 1016.500000 272.350000 1049.500000 273.650000 ;
      RECT 1007.500000 272.350000 1008.500000 273.650000 ;
      RECT 966.500000 272.350000 999.500000 273.650000 ;
      RECT 957.500000 272.350000 958.500000 273.650000 ;
      RECT 916.500000 272.350000 949.500000 273.650000 ;
      RECT 907.500000 272.350000 908.500000 273.650000 ;
      RECT 866.500000 272.350000 899.500000 273.650000 ;
      RECT 857.500000 272.350000 858.500000 273.650000 ;
      RECT 816.500000 272.350000 849.500000 273.650000 ;
      RECT 807.500000 272.350000 808.500000 273.650000 ;
      RECT 766.500000 272.350000 799.500000 273.650000 ;
      RECT 757.500000 272.350000 758.500000 273.650000 ;
      RECT 716.500000 272.350000 749.500000 273.650000 ;
      RECT 707.500000 272.350000 708.500000 273.650000 ;
      RECT 666.500000 272.350000 699.500000 273.650000 ;
      RECT 657.500000 272.350000 658.500000 273.650000 ;
      RECT 616.500000 272.350000 649.500000 273.650000 ;
      RECT 607.500000 272.350000 608.500000 273.650000 ;
      RECT 566.500000 272.350000 599.500000 273.650000 ;
      RECT 557.500000 272.350000 558.500000 273.650000 ;
      RECT 516.500000 272.350000 549.500000 273.650000 ;
      RECT 507.500000 272.350000 508.500000 273.650000 ;
      RECT 466.500000 272.350000 499.500000 273.650000 ;
      RECT 457.500000 272.350000 458.500000 273.650000 ;
      RECT 416.500000 272.350000 449.500000 273.650000 ;
      RECT 407.500000 272.350000 408.500000 273.650000 ;
      RECT 366.500000 272.350000 399.500000 273.650000 ;
      RECT 357.500000 272.350000 358.500000 273.650000 ;
      RECT 316.500000 272.350000 349.500000 273.650000 ;
      RECT 307.500000 272.350000 308.500000 273.650000 ;
      RECT 266.500000 272.350000 299.500000 273.650000 ;
      RECT 257.500000 272.350000 258.500000 273.650000 ;
      RECT 216.500000 272.350000 249.500000 273.650000 ;
      RECT 207.500000 272.350000 208.500000 273.650000 ;
      RECT 166.500000 272.350000 199.500000 273.650000 ;
      RECT 157.500000 272.350000 158.500000 273.650000 ;
      RECT 116.500000 272.350000 149.500000 273.650000 ;
      RECT 107.500000 272.350000 108.500000 273.650000 ;
      RECT 66.500000 272.350000 99.500000 273.650000 ;
      RECT 57.500000 272.350000 58.500000 273.650000 ;
      RECT 29.500000 272.350000 49.500000 273.650000 ;
      RECT 15.500000 272.350000 16.500000 273.650000 ;
      RECT 0.000000 272.350000 2.500000 275.650000 ;
      RECT 1169.500000 271.650000 1186.000000 272.350000 ;
      RECT 1116.500000 271.650000 1156.500000 272.350000 ;
      RECT 1066.500000 271.650000 1108.500000 272.350000 ;
      RECT 1016.500000 271.650000 1058.500000 272.350000 ;
      RECT 966.500000 271.650000 1008.500000 272.350000 ;
      RECT 916.500000 271.650000 958.500000 272.350000 ;
      RECT 866.500000 271.650000 908.500000 272.350000 ;
      RECT 816.500000 271.650000 858.500000 272.350000 ;
      RECT 766.500000 271.650000 808.500000 272.350000 ;
      RECT 716.500000 271.650000 758.500000 272.350000 ;
      RECT 666.500000 271.650000 708.500000 272.350000 ;
      RECT 616.500000 271.650000 658.500000 272.350000 ;
      RECT 566.500000 271.650000 608.500000 272.350000 ;
      RECT 516.500000 271.650000 558.500000 272.350000 ;
      RECT 466.500000 271.650000 508.500000 272.350000 ;
      RECT 416.500000 271.650000 458.500000 272.350000 ;
      RECT 366.500000 271.650000 408.500000 272.350000 ;
      RECT 316.500000 271.650000 358.500000 272.350000 ;
      RECT 266.500000 271.650000 308.500000 272.350000 ;
      RECT 216.500000 271.650000 258.500000 272.350000 ;
      RECT 166.500000 271.650000 208.500000 272.350000 ;
      RECT 116.500000 271.650000 158.500000 272.350000 ;
      RECT 66.500000 271.650000 108.500000 272.350000 ;
      RECT 29.500000 271.650000 58.500000 272.350000 ;
      RECT 0.000000 271.650000 16.500000 272.350000 ;
      RECT 1169.500000 270.350000 1170.500000 271.650000 ;
      RECT 1116.500000 270.350000 1149.500000 271.650000 ;
      RECT 1107.500000 270.350000 1108.500000 271.650000 ;
      RECT 1066.500000 270.350000 1099.500000 271.650000 ;
      RECT 1057.500000 270.350000 1058.500000 271.650000 ;
      RECT 1016.500000 270.350000 1049.500000 271.650000 ;
      RECT 1007.500000 270.350000 1008.500000 271.650000 ;
      RECT 966.500000 270.350000 999.500000 271.650000 ;
      RECT 957.500000 270.350000 958.500000 271.650000 ;
      RECT 916.500000 270.350000 949.500000 271.650000 ;
      RECT 907.500000 270.350000 908.500000 271.650000 ;
      RECT 866.500000 270.350000 899.500000 271.650000 ;
      RECT 857.500000 270.350000 858.500000 271.650000 ;
      RECT 816.500000 270.350000 849.500000 271.650000 ;
      RECT 807.500000 270.350000 808.500000 271.650000 ;
      RECT 766.500000 270.350000 799.500000 271.650000 ;
      RECT 757.500000 270.350000 758.500000 271.650000 ;
      RECT 716.500000 270.350000 749.500000 271.650000 ;
      RECT 707.500000 270.350000 708.500000 271.650000 ;
      RECT 666.500000 270.350000 699.500000 271.650000 ;
      RECT 657.500000 270.350000 658.500000 271.650000 ;
      RECT 616.500000 270.350000 649.500000 271.650000 ;
      RECT 607.500000 270.350000 608.500000 271.650000 ;
      RECT 566.500000 270.350000 599.500000 271.650000 ;
      RECT 557.500000 270.350000 558.500000 271.650000 ;
      RECT 516.500000 270.350000 549.500000 271.650000 ;
      RECT 507.500000 270.350000 508.500000 271.650000 ;
      RECT 466.500000 270.350000 499.500000 271.650000 ;
      RECT 457.500000 270.350000 458.500000 271.650000 ;
      RECT 416.500000 270.350000 449.500000 271.650000 ;
      RECT 407.500000 270.350000 408.500000 271.650000 ;
      RECT 366.500000 270.350000 399.500000 271.650000 ;
      RECT 357.500000 270.350000 358.500000 271.650000 ;
      RECT 316.500000 270.350000 349.500000 271.650000 ;
      RECT 307.500000 270.350000 308.500000 271.650000 ;
      RECT 266.500000 270.350000 299.500000 271.650000 ;
      RECT 257.500000 270.350000 258.500000 271.650000 ;
      RECT 216.500000 270.350000 249.500000 271.650000 ;
      RECT 207.500000 270.350000 208.500000 271.650000 ;
      RECT 166.500000 270.350000 199.500000 271.650000 ;
      RECT 157.500000 270.350000 158.500000 271.650000 ;
      RECT 116.500000 270.350000 149.500000 271.650000 ;
      RECT 107.500000 270.350000 108.500000 271.650000 ;
      RECT 66.500000 270.350000 99.500000 271.650000 ;
      RECT 57.500000 270.350000 58.500000 271.650000 ;
      RECT 29.500000 270.350000 49.500000 271.650000 ;
      RECT 15.500000 270.350000 16.500000 271.650000 ;
      RECT 1157.500000 269.650000 1170.500000 270.350000 ;
      RECT 1107.500000 269.650000 1149.500000 270.350000 ;
      RECT 1057.500000 269.650000 1099.500000 270.350000 ;
      RECT 1007.500000 269.650000 1049.500000 270.350000 ;
      RECT 957.500000 269.650000 999.500000 270.350000 ;
      RECT 907.500000 269.650000 949.500000 270.350000 ;
      RECT 857.500000 269.650000 899.500000 270.350000 ;
      RECT 807.500000 269.650000 849.500000 270.350000 ;
      RECT 757.500000 269.650000 799.500000 270.350000 ;
      RECT 707.500000 269.650000 749.500000 270.350000 ;
      RECT 657.500000 269.650000 699.500000 270.350000 ;
      RECT 607.500000 269.650000 649.500000 270.350000 ;
      RECT 557.500000 269.650000 599.500000 270.350000 ;
      RECT 507.500000 269.650000 549.500000 270.350000 ;
      RECT 457.500000 269.650000 499.500000 270.350000 ;
      RECT 407.500000 269.650000 449.500000 270.350000 ;
      RECT 357.500000 269.650000 399.500000 270.350000 ;
      RECT 307.500000 269.650000 349.500000 270.350000 ;
      RECT 257.500000 269.650000 299.500000 270.350000 ;
      RECT 207.500000 269.650000 249.500000 270.350000 ;
      RECT 157.500000 269.650000 199.500000 270.350000 ;
      RECT 107.500000 269.650000 149.500000 270.350000 ;
      RECT 57.500000 269.650000 99.500000 270.350000 ;
      RECT 15.500000 269.650000 49.500000 270.350000 ;
      RECT 1183.500000 268.350000 1186.000000 271.650000 ;
      RECT 1169.500000 268.350000 1170.500000 269.650000 ;
      RECT 1116.500000 268.350000 1149.500000 269.650000 ;
      RECT 1107.500000 268.350000 1108.500000 269.650000 ;
      RECT 1066.500000 268.350000 1099.500000 269.650000 ;
      RECT 1057.500000 268.350000 1058.500000 269.650000 ;
      RECT 1016.500000 268.350000 1049.500000 269.650000 ;
      RECT 1007.500000 268.350000 1008.500000 269.650000 ;
      RECT 966.500000 268.350000 999.500000 269.650000 ;
      RECT 957.500000 268.350000 958.500000 269.650000 ;
      RECT 916.500000 268.350000 949.500000 269.650000 ;
      RECT 907.500000 268.350000 908.500000 269.650000 ;
      RECT 866.500000 268.350000 899.500000 269.650000 ;
      RECT 857.500000 268.350000 858.500000 269.650000 ;
      RECT 816.500000 268.350000 849.500000 269.650000 ;
      RECT 807.500000 268.350000 808.500000 269.650000 ;
      RECT 766.500000 268.350000 799.500000 269.650000 ;
      RECT 757.500000 268.350000 758.500000 269.650000 ;
      RECT 716.500000 268.350000 749.500000 269.650000 ;
      RECT 707.500000 268.350000 708.500000 269.650000 ;
      RECT 666.500000 268.350000 699.500000 269.650000 ;
      RECT 657.500000 268.350000 658.500000 269.650000 ;
      RECT 616.500000 268.350000 649.500000 269.650000 ;
      RECT 607.500000 268.350000 608.500000 269.650000 ;
      RECT 566.500000 268.350000 599.500000 269.650000 ;
      RECT 557.500000 268.350000 558.500000 269.650000 ;
      RECT 516.500000 268.350000 549.500000 269.650000 ;
      RECT 507.500000 268.350000 508.500000 269.650000 ;
      RECT 466.500000 268.350000 499.500000 269.650000 ;
      RECT 457.500000 268.350000 458.500000 269.650000 ;
      RECT 416.500000 268.350000 449.500000 269.650000 ;
      RECT 407.500000 268.350000 408.500000 269.650000 ;
      RECT 366.500000 268.350000 399.500000 269.650000 ;
      RECT 357.500000 268.350000 358.500000 269.650000 ;
      RECT 316.500000 268.350000 349.500000 269.650000 ;
      RECT 307.500000 268.350000 308.500000 269.650000 ;
      RECT 266.500000 268.350000 299.500000 269.650000 ;
      RECT 257.500000 268.350000 258.500000 269.650000 ;
      RECT 216.500000 268.350000 249.500000 269.650000 ;
      RECT 207.500000 268.350000 208.500000 269.650000 ;
      RECT 166.500000 268.350000 199.500000 269.650000 ;
      RECT 157.500000 268.350000 158.500000 269.650000 ;
      RECT 116.500000 268.350000 149.500000 269.650000 ;
      RECT 107.500000 268.350000 108.500000 269.650000 ;
      RECT 66.500000 268.350000 99.500000 269.650000 ;
      RECT 57.500000 268.350000 58.500000 269.650000 ;
      RECT 29.500000 268.350000 49.500000 269.650000 ;
      RECT 15.500000 268.350000 16.500000 269.650000 ;
      RECT 0.000000 268.350000 2.500000 271.650000 ;
      RECT 1169.500000 267.650000 1186.000000 268.350000 ;
      RECT 1116.500000 267.650000 1156.500000 268.350000 ;
      RECT 1066.500000 267.650000 1108.500000 268.350000 ;
      RECT 1016.500000 267.650000 1058.500000 268.350000 ;
      RECT 966.500000 267.650000 1008.500000 268.350000 ;
      RECT 916.500000 267.650000 958.500000 268.350000 ;
      RECT 866.500000 267.650000 908.500000 268.350000 ;
      RECT 816.500000 267.650000 858.500000 268.350000 ;
      RECT 766.500000 267.650000 808.500000 268.350000 ;
      RECT 716.500000 267.650000 758.500000 268.350000 ;
      RECT 666.500000 267.650000 708.500000 268.350000 ;
      RECT 616.500000 267.650000 658.500000 268.350000 ;
      RECT 566.500000 267.650000 608.500000 268.350000 ;
      RECT 516.500000 267.650000 558.500000 268.350000 ;
      RECT 466.500000 267.650000 508.500000 268.350000 ;
      RECT 416.500000 267.650000 458.500000 268.350000 ;
      RECT 366.500000 267.650000 408.500000 268.350000 ;
      RECT 316.500000 267.650000 358.500000 268.350000 ;
      RECT 266.500000 267.650000 308.500000 268.350000 ;
      RECT 216.500000 267.650000 258.500000 268.350000 ;
      RECT 166.500000 267.650000 208.500000 268.350000 ;
      RECT 116.500000 267.650000 158.500000 268.350000 ;
      RECT 66.500000 267.650000 108.500000 268.350000 ;
      RECT 29.500000 267.650000 58.500000 268.350000 ;
      RECT 0.000000 267.650000 16.500000 268.350000 ;
      RECT 1169.500000 266.350000 1170.500000 267.650000 ;
      RECT 1116.500000 266.350000 1149.500000 267.650000 ;
      RECT 1107.500000 266.350000 1108.500000 267.650000 ;
      RECT 1066.500000 266.350000 1099.500000 267.650000 ;
      RECT 1057.500000 266.350000 1058.500000 267.650000 ;
      RECT 1016.500000 266.350000 1049.500000 267.650000 ;
      RECT 1007.500000 266.350000 1008.500000 267.650000 ;
      RECT 966.500000 266.350000 999.500000 267.650000 ;
      RECT 957.500000 266.350000 958.500000 267.650000 ;
      RECT 916.500000 266.350000 949.500000 267.650000 ;
      RECT 907.500000 266.350000 908.500000 267.650000 ;
      RECT 866.500000 266.350000 899.500000 267.650000 ;
      RECT 857.500000 266.350000 858.500000 267.650000 ;
      RECT 816.500000 266.350000 849.500000 267.650000 ;
      RECT 807.500000 266.350000 808.500000 267.650000 ;
      RECT 766.500000 266.350000 799.500000 267.650000 ;
      RECT 757.500000 266.350000 758.500000 267.650000 ;
      RECT 716.500000 266.350000 749.500000 267.650000 ;
      RECT 707.500000 266.350000 708.500000 267.650000 ;
      RECT 666.500000 266.350000 699.500000 267.650000 ;
      RECT 657.500000 266.350000 658.500000 267.650000 ;
      RECT 616.500000 266.350000 649.500000 267.650000 ;
      RECT 607.500000 266.350000 608.500000 267.650000 ;
      RECT 566.500000 266.350000 599.500000 267.650000 ;
      RECT 557.500000 266.350000 558.500000 267.650000 ;
      RECT 516.500000 266.350000 549.500000 267.650000 ;
      RECT 507.500000 266.350000 508.500000 267.650000 ;
      RECT 466.500000 266.350000 499.500000 267.650000 ;
      RECT 457.500000 266.350000 458.500000 267.650000 ;
      RECT 416.500000 266.350000 449.500000 267.650000 ;
      RECT 407.500000 266.350000 408.500000 267.650000 ;
      RECT 366.500000 266.350000 399.500000 267.650000 ;
      RECT 357.500000 266.350000 358.500000 267.650000 ;
      RECT 316.500000 266.350000 349.500000 267.650000 ;
      RECT 307.500000 266.350000 308.500000 267.650000 ;
      RECT 266.500000 266.350000 299.500000 267.650000 ;
      RECT 257.500000 266.350000 258.500000 267.650000 ;
      RECT 216.500000 266.350000 249.500000 267.650000 ;
      RECT 207.500000 266.350000 208.500000 267.650000 ;
      RECT 166.500000 266.350000 199.500000 267.650000 ;
      RECT 157.500000 266.350000 158.500000 267.650000 ;
      RECT 116.500000 266.350000 149.500000 267.650000 ;
      RECT 107.500000 266.350000 108.500000 267.650000 ;
      RECT 66.500000 266.350000 99.500000 267.650000 ;
      RECT 57.500000 266.350000 58.500000 267.650000 ;
      RECT 29.500000 266.350000 49.500000 267.650000 ;
      RECT 15.500000 266.350000 16.500000 267.650000 ;
      RECT 1157.500000 265.650000 1170.500000 266.350000 ;
      RECT 1107.500000 265.650000 1149.500000 266.350000 ;
      RECT 1057.500000 265.650000 1099.500000 266.350000 ;
      RECT 1007.500000 265.650000 1049.500000 266.350000 ;
      RECT 957.500000 265.650000 999.500000 266.350000 ;
      RECT 907.500000 265.650000 949.500000 266.350000 ;
      RECT 857.500000 265.650000 899.500000 266.350000 ;
      RECT 807.500000 265.650000 849.500000 266.350000 ;
      RECT 757.500000 265.650000 799.500000 266.350000 ;
      RECT 707.500000 265.650000 749.500000 266.350000 ;
      RECT 657.500000 265.650000 699.500000 266.350000 ;
      RECT 607.500000 265.650000 649.500000 266.350000 ;
      RECT 557.500000 265.650000 599.500000 266.350000 ;
      RECT 507.500000 265.650000 549.500000 266.350000 ;
      RECT 457.500000 265.650000 499.500000 266.350000 ;
      RECT 407.500000 265.650000 449.500000 266.350000 ;
      RECT 357.500000 265.650000 399.500000 266.350000 ;
      RECT 307.500000 265.650000 349.500000 266.350000 ;
      RECT 257.500000 265.650000 299.500000 266.350000 ;
      RECT 207.500000 265.650000 249.500000 266.350000 ;
      RECT 157.500000 265.650000 199.500000 266.350000 ;
      RECT 107.500000 265.650000 149.500000 266.350000 ;
      RECT 57.500000 265.650000 99.500000 266.350000 ;
      RECT 15.500000 265.650000 49.500000 266.350000 ;
      RECT 1183.500000 264.350000 1186.000000 267.650000 ;
      RECT 1169.500000 264.350000 1170.500000 265.650000 ;
      RECT 1116.500000 264.350000 1149.500000 265.650000 ;
      RECT 1107.500000 264.350000 1108.500000 265.650000 ;
      RECT 1066.500000 264.350000 1099.500000 265.650000 ;
      RECT 1057.500000 264.350000 1058.500000 265.650000 ;
      RECT 1016.500000 264.350000 1049.500000 265.650000 ;
      RECT 1007.500000 264.350000 1008.500000 265.650000 ;
      RECT 966.500000 264.350000 999.500000 265.650000 ;
      RECT 957.500000 264.350000 958.500000 265.650000 ;
      RECT 916.500000 264.350000 949.500000 265.650000 ;
      RECT 907.500000 264.350000 908.500000 265.650000 ;
      RECT 866.500000 264.350000 899.500000 265.650000 ;
      RECT 857.500000 264.350000 858.500000 265.650000 ;
      RECT 816.500000 264.350000 849.500000 265.650000 ;
      RECT 807.500000 264.350000 808.500000 265.650000 ;
      RECT 766.500000 264.350000 799.500000 265.650000 ;
      RECT 757.500000 264.350000 758.500000 265.650000 ;
      RECT 716.500000 264.350000 749.500000 265.650000 ;
      RECT 707.500000 264.350000 708.500000 265.650000 ;
      RECT 666.500000 264.350000 699.500000 265.650000 ;
      RECT 657.500000 264.350000 658.500000 265.650000 ;
      RECT 616.500000 264.350000 649.500000 265.650000 ;
      RECT 607.500000 264.350000 608.500000 265.650000 ;
      RECT 566.500000 264.350000 599.500000 265.650000 ;
      RECT 557.500000 264.350000 558.500000 265.650000 ;
      RECT 516.500000 264.350000 549.500000 265.650000 ;
      RECT 507.500000 264.350000 508.500000 265.650000 ;
      RECT 466.500000 264.350000 499.500000 265.650000 ;
      RECT 457.500000 264.350000 458.500000 265.650000 ;
      RECT 416.500000 264.350000 449.500000 265.650000 ;
      RECT 407.500000 264.350000 408.500000 265.650000 ;
      RECT 366.500000 264.350000 399.500000 265.650000 ;
      RECT 357.500000 264.350000 358.500000 265.650000 ;
      RECT 316.500000 264.350000 349.500000 265.650000 ;
      RECT 307.500000 264.350000 308.500000 265.650000 ;
      RECT 266.500000 264.350000 299.500000 265.650000 ;
      RECT 257.500000 264.350000 258.500000 265.650000 ;
      RECT 216.500000 264.350000 249.500000 265.650000 ;
      RECT 207.500000 264.350000 208.500000 265.650000 ;
      RECT 166.500000 264.350000 199.500000 265.650000 ;
      RECT 157.500000 264.350000 158.500000 265.650000 ;
      RECT 116.500000 264.350000 149.500000 265.650000 ;
      RECT 107.500000 264.350000 108.500000 265.650000 ;
      RECT 66.500000 264.350000 99.500000 265.650000 ;
      RECT 57.500000 264.350000 58.500000 265.650000 ;
      RECT 29.500000 264.350000 49.500000 265.650000 ;
      RECT 15.500000 264.350000 16.500000 265.650000 ;
      RECT 0.000000 264.350000 2.500000 267.650000 ;
      RECT 1169.500000 263.650000 1186.000000 264.350000 ;
      RECT 1116.500000 263.650000 1156.500000 264.350000 ;
      RECT 1066.500000 263.650000 1108.500000 264.350000 ;
      RECT 1016.500000 263.650000 1058.500000 264.350000 ;
      RECT 966.500000 263.650000 1008.500000 264.350000 ;
      RECT 916.500000 263.650000 958.500000 264.350000 ;
      RECT 866.500000 263.650000 908.500000 264.350000 ;
      RECT 816.500000 263.650000 858.500000 264.350000 ;
      RECT 766.500000 263.650000 808.500000 264.350000 ;
      RECT 716.500000 263.650000 758.500000 264.350000 ;
      RECT 666.500000 263.650000 708.500000 264.350000 ;
      RECT 616.500000 263.650000 658.500000 264.350000 ;
      RECT 566.500000 263.650000 608.500000 264.350000 ;
      RECT 516.500000 263.650000 558.500000 264.350000 ;
      RECT 466.500000 263.650000 508.500000 264.350000 ;
      RECT 416.500000 263.650000 458.500000 264.350000 ;
      RECT 366.500000 263.650000 408.500000 264.350000 ;
      RECT 316.500000 263.650000 358.500000 264.350000 ;
      RECT 266.500000 263.650000 308.500000 264.350000 ;
      RECT 216.500000 263.650000 258.500000 264.350000 ;
      RECT 166.500000 263.650000 208.500000 264.350000 ;
      RECT 116.500000 263.650000 158.500000 264.350000 ;
      RECT 66.500000 263.650000 108.500000 264.350000 ;
      RECT 29.500000 263.650000 58.500000 264.350000 ;
      RECT 0.000000 263.650000 16.500000 264.350000 ;
      RECT 1169.500000 262.350000 1170.500000 263.650000 ;
      RECT 1116.500000 262.350000 1149.500000 263.650000 ;
      RECT 1107.500000 262.350000 1108.500000 263.650000 ;
      RECT 1066.500000 262.350000 1099.500000 263.650000 ;
      RECT 1057.500000 262.350000 1058.500000 263.650000 ;
      RECT 1016.500000 262.350000 1049.500000 263.650000 ;
      RECT 1007.500000 262.350000 1008.500000 263.650000 ;
      RECT 966.500000 262.350000 999.500000 263.650000 ;
      RECT 957.500000 262.350000 958.500000 263.650000 ;
      RECT 916.500000 262.350000 949.500000 263.650000 ;
      RECT 907.500000 262.350000 908.500000 263.650000 ;
      RECT 866.500000 262.350000 899.500000 263.650000 ;
      RECT 857.500000 262.350000 858.500000 263.650000 ;
      RECT 816.500000 262.350000 849.500000 263.650000 ;
      RECT 807.500000 262.350000 808.500000 263.650000 ;
      RECT 766.500000 262.350000 799.500000 263.650000 ;
      RECT 757.500000 262.350000 758.500000 263.650000 ;
      RECT 716.500000 262.350000 749.500000 263.650000 ;
      RECT 707.500000 262.350000 708.500000 263.650000 ;
      RECT 666.500000 262.350000 699.500000 263.650000 ;
      RECT 657.500000 262.350000 658.500000 263.650000 ;
      RECT 616.500000 262.350000 649.500000 263.650000 ;
      RECT 607.500000 262.350000 608.500000 263.650000 ;
      RECT 566.500000 262.350000 599.500000 263.650000 ;
      RECT 557.500000 262.350000 558.500000 263.650000 ;
      RECT 516.500000 262.350000 549.500000 263.650000 ;
      RECT 507.500000 262.350000 508.500000 263.650000 ;
      RECT 466.500000 262.350000 499.500000 263.650000 ;
      RECT 457.500000 262.350000 458.500000 263.650000 ;
      RECT 416.500000 262.350000 449.500000 263.650000 ;
      RECT 407.500000 262.350000 408.500000 263.650000 ;
      RECT 366.500000 262.350000 399.500000 263.650000 ;
      RECT 357.500000 262.350000 358.500000 263.650000 ;
      RECT 316.500000 262.350000 349.500000 263.650000 ;
      RECT 307.500000 262.350000 308.500000 263.650000 ;
      RECT 266.500000 262.350000 299.500000 263.650000 ;
      RECT 257.500000 262.350000 258.500000 263.650000 ;
      RECT 216.500000 262.350000 249.500000 263.650000 ;
      RECT 207.500000 262.350000 208.500000 263.650000 ;
      RECT 166.500000 262.350000 199.500000 263.650000 ;
      RECT 157.500000 262.350000 158.500000 263.650000 ;
      RECT 116.500000 262.350000 149.500000 263.650000 ;
      RECT 107.500000 262.350000 108.500000 263.650000 ;
      RECT 66.500000 262.350000 99.500000 263.650000 ;
      RECT 57.500000 262.350000 58.500000 263.650000 ;
      RECT 29.500000 262.350000 49.500000 263.650000 ;
      RECT 15.500000 262.350000 16.500000 263.650000 ;
      RECT 1157.500000 261.650000 1170.500000 262.350000 ;
      RECT 1107.500000 261.650000 1149.500000 262.350000 ;
      RECT 1057.500000 261.650000 1099.500000 262.350000 ;
      RECT 1007.500000 261.650000 1049.500000 262.350000 ;
      RECT 957.500000 261.650000 999.500000 262.350000 ;
      RECT 907.500000 261.650000 949.500000 262.350000 ;
      RECT 857.500000 261.650000 899.500000 262.350000 ;
      RECT 807.500000 261.650000 849.500000 262.350000 ;
      RECT 757.500000 261.650000 799.500000 262.350000 ;
      RECT 707.500000 261.650000 749.500000 262.350000 ;
      RECT 657.500000 261.650000 699.500000 262.350000 ;
      RECT 607.500000 261.650000 649.500000 262.350000 ;
      RECT 557.500000 261.650000 599.500000 262.350000 ;
      RECT 507.500000 261.650000 549.500000 262.350000 ;
      RECT 457.500000 261.650000 499.500000 262.350000 ;
      RECT 407.500000 261.650000 449.500000 262.350000 ;
      RECT 357.500000 261.650000 399.500000 262.350000 ;
      RECT 307.500000 261.650000 349.500000 262.350000 ;
      RECT 257.500000 261.650000 299.500000 262.350000 ;
      RECT 207.500000 261.650000 249.500000 262.350000 ;
      RECT 157.500000 261.650000 199.500000 262.350000 ;
      RECT 107.500000 261.650000 149.500000 262.350000 ;
      RECT 57.500000 261.650000 99.500000 262.350000 ;
      RECT 15.500000 261.650000 49.500000 262.350000 ;
      RECT 1183.500000 260.350000 1186.000000 263.650000 ;
      RECT 1169.500000 260.350000 1170.500000 261.650000 ;
      RECT 1116.500000 260.350000 1149.500000 261.650000 ;
      RECT 1107.500000 260.350000 1108.500000 261.650000 ;
      RECT 1066.500000 260.350000 1099.500000 261.650000 ;
      RECT 1057.500000 260.350000 1058.500000 261.650000 ;
      RECT 1016.500000 260.350000 1049.500000 261.650000 ;
      RECT 1007.500000 260.350000 1008.500000 261.650000 ;
      RECT 966.500000 260.350000 999.500000 261.650000 ;
      RECT 957.500000 260.350000 958.500000 261.650000 ;
      RECT 916.500000 260.350000 949.500000 261.650000 ;
      RECT 907.500000 260.350000 908.500000 261.650000 ;
      RECT 866.500000 260.350000 899.500000 261.650000 ;
      RECT 857.500000 260.350000 858.500000 261.650000 ;
      RECT 816.500000 260.350000 849.500000 261.650000 ;
      RECT 807.500000 260.350000 808.500000 261.650000 ;
      RECT 766.500000 260.350000 799.500000 261.650000 ;
      RECT 757.500000 260.350000 758.500000 261.650000 ;
      RECT 716.500000 260.350000 749.500000 261.650000 ;
      RECT 707.500000 260.350000 708.500000 261.650000 ;
      RECT 666.500000 260.350000 699.500000 261.650000 ;
      RECT 657.500000 260.350000 658.500000 261.650000 ;
      RECT 616.500000 260.350000 649.500000 261.650000 ;
      RECT 607.500000 260.350000 608.500000 261.650000 ;
      RECT 566.500000 260.350000 599.500000 261.650000 ;
      RECT 557.500000 260.350000 558.500000 261.650000 ;
      RECT 516.500000 260.350000 549.500000 261.650000 ;
      RECT 507.500000 260.350000 508.500000 261.650000 ;
      RECT 466.500000 260.350000 499.500000 261.650000 ;
      RECT 457.500000 260.350000 458.500000 261.650000 ;
      RECT 416.500000 260.350000 449.500000 261.650000 ;
      RECT 407.500000 260.350000 408.500000 261.650000 ;
      RECT 366.500000 260.350000 399.500000 261.650000 ;
      RECT 357.500000 260.350000 358.500000 261.650000 ;
      RECT 316.500000 260.350000 349.500000 261.650000 ;
      RECT 307.500000 260.350000 308.500000 261.650000 ;
      RECT 266.500000 260.350000 299.500000 261.650000 ;
      RECT 257.500000 260.350000 258.500000 261.650000 ;
      RECT 216.500000 260.350000 249.500000 261.650000 ;
      RECT 207.500000 260.350000 208.500000 261.650000 ;
      RECT 166.500000 260.350000 199.500000 261.650000 ;
      RECT 157.500000 260.350000 158.500000 261.650000 ;
      RECT 116.500000 260.350000 149.500000 261.650000 ;
      RECT 107.500000 260.350000 108.500000 261.650000 ;
      RECT 66.500000 260.350000 99.500000 261.650000 ;
      RECT 57.500000 260.350000 58.500000 261.650000 ;
      RECT 29.500000 260.350000 49.500000 261.650000 ;
      RECT 15.500000 260.350000 16.500000 261.650000 ;
      RECT 0.000000 260.350000 2.500000 263.650000 ;
      RECT 1169.500000 259.650000 1186.000000 260.350000 ;
      RECT 1116.500000 259.650000 1156.500000 260.350000 ;
      RECT 1169.500000 258.350000 1170.500000 259.650000 ;
      RECT 1116.500000 258.350000 1149.500000 259.650000 ;
      RECT 1066.500000 258.350000 1108.500000 260.350000 ;
      RECT 1016.500000 258.350000 1058.500000 260.350000 ;
      RECT 966.500000 258.350000 1008.500000 260.350000 ;
      RECT 916.500000 258.350000 958.500000 260.350000 ;
      RECT 866.500000 258.350000 908.500000 260.350000 ;
      RECT 816.500000 258.350000 858.500000 260.350000 ;
      RECT 766.500000 258.350000 808.500000 260.350000 ;
      RECT 716.500000 258.350000 758.500000 260.350000 ;
      RECT 666.500000 258.350000 708.500000 260.350000 ;
      RECT 616.500000 258.350000 658.500000 260.350000 ;
      RECT 566.500000 258.350000 608.500000 260.350000 ;
      RECT 516.500000 258.350000 558.500000 260.350000 ;
      RECT 466.500000 258.350000 508.500000 260.350000 ;
      RECT 416.500000 258.350000 458.500000 260.350000 ;
      RECT 366.500000 258.350000 408.500000 260.350000 ;
      RECT 316.500000 258.350000 358.500000 260.350000 ;
      RECT 266.500000 258.350000 308.500000 260.350000 ;
      RECT 216.500000 258.350000 258.500000 260.350000 ;
      RECT 166.500000 258.350000 208.500000 260.350000 ;
      RECT 116.500000 258.350000 158.500000 260.350000 ;
      RECT 66.500000 258.350000 108.500000 260.350000 ;
      RECT 29.500000 258.350000 58.500000 260.350000 ;
      RECT 0.000000 258.350000 16.500000 260.350000 ;
      RECT 1157.500000 257.650000 1170.500000 258.350000 ;
      RECT 1183.500000 256.350000 1186.000000 259.650000 ;
      RECT 1169.500000 256.350000 1170.500000 257.650000 ;
      RECT 0.000000 256.350000 1149.500000 258.350000 ;
      RECT 1169.500000 255.650000 1186.000000 256.350000 ;
      RECT 1169.500000 254.350000 1170.500000 255.650000 ;
      RECT 0.000000 254.350000 1156.500000 256.350000 ;
      RECT 0.000000 253.650000 1170.500000 254.350000 ;
      RECT 1183.500000 252.350000 1186.000000 255.650000 ;
      RECT 1169.500000 252.350000 1170.500000 253.650000 ;
      RECT 1169.500000 251.650000 1186.000000 252.350000 ;
      RECT 1169.500000 250.350000 1170.500000 251.650000 ;
      RECT 0.000000 250.350000 1156.500000 253.650000 ;
      RECT 0.000000 249.650000 1170.500000 250.350000 ;
      RECT 1183.500000 248.350000 1186.000000 251.650000 ;
      RECT 1169.500000 248.350000 1170.500000 249.650000 ;
      RECT 1169.500000 247.650000 1186.000000 248.350000 ;
      RECT 1169.500000 246.350000 1170.500000 247.650000 ;
      RECT 0.000000 246.350000 1156.500000 249.650000 ;
      RECT 0.000000 245.650000 1170.500000 246.350000 ;
      RECT 1183.500000 244.350000 1186.000000 247.650000 ;
      RECT 1169.500000 244.350000 1170.500000 245.650000 ;
      RECT 1169.500000 243.650000 1186.000000 244.350000 ;
      RECT 1169.500000 242.350000 1170.500000 243.650000 ;
      RECT 0.000000 242.350000 1156.500000 245.650000 ;
      RECT 0.000000 241.650000 1170.500000 242.350000 ;
      RECT 1183.500000 240.350000 1186.000000 243.650000 ;
      RECT 1169.500000 240.350000 1170.500000 241.650000 ;
      RECT 1169.500000 239.650000 1186.000000 240.350000 ;
      RECT 1169.500000 238.350000 1170.500000 239.650000 ;
      RECT 0.000000 238.350000 1156.500000 241.650000 ;
      RECT 0.000000 237.650000 1170.500000 238.350000 ;
      RECT 1183.500000 236.350000 1186.000000 239.650000 ;
      RECT 1169.500000 236.350000 1170.500000 237.650000 ;
      RECT 1169.500000 235.650000 1186.000000 236.350000 ;
      RECT 1169.500000 234.350000 1170.500000 235.650000 ;
      RECT 0.000000 234.350000 1156.500000 237.650000 ;
      RECT 0.000000 233.650000 1170.500000 234.350000 ;
      RECT 1183.500000 232.350000 1186.000000 235.650000 ;
      RECT 1169.500000 232.350000 1170.500000 233.650000 ;
      RECT 1169.500000 231.650000 1186.000000 232.350000 ;
      RECT 1169.500000 230.350000 1170.500000 231.650000 ;
      RECT 0.000000 230.350000 1156.500000 233.650000 ;
      RECT 0.000000 229.650000 1170.500000 230.350000 ;
      RECT 1183.500000 228.350000 1186.000000 231.650000 ;
      RECT 1169.500000 228.350000 1170.500000 229.650000 ;
      RECT 1169.500000 227.650000 1186.000000 228.350000 ;
      RECT 1169.500000 226.350000 1170.500000 227.650000 ;
      RECT 0.000000 226.350000 1156.500000 229.650000 ;
      RECT 0.000000 225.650000 1170.500000 226.350000 ;
      RECT 1183.500000 224.350000 1186.000000 227.650000 ;
      RECT 1169.500000 224.350000 1170.500000 225.650000 ;
      RECT 1169.500000 223.650000 1186.000000 224.350000 ;
      RECT 0.000000 223.170000 1156.500000 225.650000 ;
      RECT 1183.500000 223.165000 1186.000000 223.650000 ;
      RECT 1169.500000 222.350000 1170.500000 223.650000 ;
      RECT 2.020000 222.350000 1156.500000 223.170000 ;
      RECT 2.020000 221.650000 1170.500000 222.350000 ;
      RECT 1183.500000 220.350000 1183.980000 223.165000 ;
      RECT 1169.500000 220.350000 1170.500000 221.650000 ;
      RECT 2.020000 220.070000 1156.500000 221.650000 ;
      RECT 1169.500000 220.065000 1183.980000 220.350000 ;
      RECT 1169.500000 219.650000 1186.000000 220.065000 ;
      RECT 1169.500000 218.350000 1170.500000 219.650000 ;
      RECT 0.000000 218.350000 1156.500000 220.070000 ;
      RECT 0.000000 217.650000 1170.500000 218.350000 ;
      RECT 1183.500000 217.485000 1186.000000 219.650000 ;
      RECT 1183.500000 216.350000 1183.980000 217.485000 ;
      RECT 1169.500000 216.350000 1170.500000 217.650000 ;
      RECT 1169.500000 215.650000 1183.980000 216.350000 ;
      RECT 1183.500000 214.385000 1183.980000 215.650000 ;
      RECT 1169.500000 214.350000 1170.500000 215.650000 ;
      RECT 0.000000 214.350000 1156.500000 217.650000 ;
      RECT 0.000000 213.650000 1170.500000 214.350000 ;
      RECT 1183.500000 213.525000 1186.000000 214.385000 ;
      RECT 0.000000 212.575000 1156.500000 213.650000 ;
      RECT 1183.500000 212.350000 1183.980000 213.525000 ;
      RECT 1169.500000 212.350000 1170.500000 213.650000 ;
      RECT 1169.500000 211.650000 1183.980000 212.350000 ;
      RECT 1183.500000 210.425000 1183.980000 211.650000 ;
      RECT 1169.500000 210.350000 1170.500000 211.650000 ;
      RECT 2.020000 210.350000 1156.500000 212.575000 ;
      RECT 2.020000 209.650000 1170.500000 210.350000 ;
      RECT 2.020000 209.475000 1156.500000 209.650000 ;
      RECT 0.000000 208.615000 1156.500000 209.475000 ;
      RECT 1183.500000 208.350000 1186.000000 210.425000 ;
      RECT 1169.500000 208.350000 1170.500000 209.650000 ;
      RECT 1169.500000 207.650000 1186.000000 208.350000 ;
      RECT 1169.500000 206.350000 1170.500000 207.650000 ;
      RECT 2.020000 206.350000 1156.500000 208.615000 ;
      RECT 2.020000 205.650000 1170.500000 206.350000 ;
      RECT 2.020000 205.515000 1156.500000 205.650000 ;
      RECT 1183.500000 204.350000 1186.000000 207.650000 ;
      RECT 1169.500000 204.350000 1170.500000 205.650000 ;
      RECT 1169.500000 203.650000 1186.000000 204.350000 ;
      RECT 0.000000 202.935000 1156.500000 205.515000 ;
      RECT 1183.500000 202.930000 1186.000000 203.650000 ;
      RECT 1169.500000 202.350000 1170.500000 203.650000 ;
      RECT 2.020000 202.350000 1156.500000 202.935000 ;
      RECT 2.020000 201.650000 1170.500000 202.350000 ;
      RECT 1183.500000 200.350000 1183.980000 202.930000 ;
      RECT 1169.500000 200.350000 1170.500000 201.650000 ;
      RECT 2.020000 199.835000 1156.500000 201.650000 ;
      RECT 1169.500000 199.830000 1183.980000 200.350000 ;
      RECT 1169.500000 199.650000 1186.000000 199.830000 ;
      RECT 1169.500000 198.350000 1170.500000 199.650000 ;
      RECT 0.000000 198.350000 1156.500000 199.835000 ;
      RECT 0.000000 197.650000 1170.500000 198.350000 ;
      RECT 1183.500000 196.350000 1186.000000 199.650000 ;
      RECT 1169.500000 196.350000 1170.500000 197.650000 ;
      RECT 1169.500000 195.650000 1186.000000 196.350000 ;
      RECT 1169.500000 194.350000 1170.500000 195.650000 ;
      RECT 0.000000 194.350000 1156.500000 197.650000 ;
      RECT 0.000000 193.650000 1170.500000 194.350000 ;
      RECT 1183.500000 192.350000 1186.000000 195.650000 ;
      RECT 1169.500000 192.350000 1170.500000 193.650000 ;
      RECT 1169.500000 191.650000 1186.000000 192.350000 ;
      RECT 1169.500000 190.350000 1170.500000 191.650000 ;
      RECT 0.000000 190.350000 1156.500000 193.650000 ;
      RECT 0.000000 189.650000 1170.500000 190.350000 ;
      RECT 1183.500000 188.350000 1186.000000 191.650000 ;
      RECT 1169.500000 188.350000 1170.500000 189.650000 ;
      RECT 1169.500000 187.650000 1186.000000 188.350000 ;
      RECT 1169.500000 186.350000 1170.500000 187.650000 ;
      RECT 0.000000 186.350000 1156.500000 189.650000 ;
      RECT 0.000000 185.650000 1170.500000 186.350000 ;
      RECT 1183.500000 184.350000 1186.000000 187.650000 ;
      RECT 1169.500000 184.350000 1170.500000 185.650000 ;
      RECT 1169.500000 183.650000 1186.000000 184.350000 ;
      RECT 1169.500000 182.350000 1170.500000 183.650000 ;
      RECT 0.000000 182.350000 1156.500000 185.650000 ;
      RECT 0.000000 181.650000 1170.500000 182.350000 ;
      RECT 1183.500000 180.350000 1186.000000 183.650000 ;
      RECT 1169.500000 180.350000 1170.500000 181.650000 ;
      RECT 1169.500000 179.650000 1186.000000 180.350000 ;
      RECT 1169.500000 178.350000 1170.500000 179.650000 ;
      RECT 0.000000 178.350000 1156.500000 181.650000 ;
      RECT 0.000000 177.650000 1170.500000 178.350000 ;
      RECT 1183.500000 176.350000 1186.000000 179.650000 ;
      RECT 1169.500000 176.350000 1170.500000 177.650000 ;
      RECT 1169.500000 175.650000 1186.000000 176.350000 ;
      RECT 1169.500000 174.350000 1170.500000 175.650000 ;
      RECT 0.000000 174.350000 1156.500000 177.650000 ;
      RECT 0.000000 173.650000 1170.500000 174.350000 ;
      RECT 1183.500000 172.350000 1186.000000 175.650000 ;
      RECT 1169.500000 172.350000 1170.500000 173.650000 ;
      RECT 1169.500000 171.650000 1186.000000 172.350000 ;
      RECT 1169.500000 170.350000 1170.500000 171.650000 ;
      RECT 0.000000 170.350000 1156.500000 173.650000 ;
      RECT 0.000000 169.650000 1170.500000 170.350000 ;
      RECT 1183.500000 168.350000 1186.000000 171.650000 ;
      RECT 1169.500000 168.350000 1170.500000 169.650000 ;
      RECT 1169.500000 167.650000 1186.000000 168.350000 ;
      RECT 1169.500000 166.350000 1170.500000 167.650000 ;
      RECT 0.000000 166.350000 1156.500000 169.650000 ;
      RECT 0.000000 165.650000 1170.500000 166.350000 ;
      RECT 1183.500000 164.350000 1186.000000 167.650000 ;
      RECT 1169.500000 164.350000 1170.500000 165.650000 ;
      RECT 1169.500000 163.650000 1186.000000 164.350000 ;
      RECT 1169.500000 162.350000 1170.500000 163.650000 ;
      RECT 0.000000 162.350000 1156.500000 165.650000 ;
      RECT 0.000000 161.650000 1170.500000 162.350000 ;
      RECT 1183.500000 160.350000 1186.000000 163.650000 ;
      RECT 1169.500000 160.350000 1170.500000 161.650000 ;
      RECT 1169.500000 159.650000 1186.000000 160.350000 ;
      RECT 1169.500000 158.350000 1170.500000 159.650000 ;
      RECT 0.000000 158.350000 1156.500000 161.650000 ;
      RECT 0.000000 157.650000 1170.500000 158.350000 ;
      RECT 1183.500000 156.350000 1186.000000 159.650000 ;
      RECT 1169.500000 156.350000 1170.500000 157.650000 ;
      RECT 1169.500000 155.650000 1186.000000 156.350000 ;
      RECT 1169.500000 154.350000 1170.500000 155.650000 ;
      RECT 0.000000 154.350000 1156.500000 157.650000 ;
      RECT 0.000000 153.650000 1170.500000 154.350000 ;
      RECT 1183.500000 152.350000 1186.000000 155.650000 ;
      RECT 1169.500000 152.350000 1170.500000 153.650000 ;
      RECT 1169.500000 151.650000 1186.000000 152.350000 ;
      RECT 1169.500000 150.350000 1170.500000 151.650000 ;
      RECT 0.000000 150.350000 1156.500000 153.650000 ;
      RECT 0.000000 149.650000 1170.500000 150.350000 ;
      RECT 1183.500000 148.350000 1186.000000 151.650000 ;
      RECT 1169.500000 148.350000 1170.500000 149.650000 ;
      RECT 1169.500000 147.650000 1186.000000 148.350000 ;
      RECT 1169.500000 146.350000 1170.500000 147.650000 ;
      RECT 0.000000 146.350000 1156.500000 149.650000 ;
      RECT 0.000000 145.650000 1170.500000 146.350000 ;
      RECT 1183.500000 144.350000 1186.000000 147.650000 ;
      RECT 1169.500000 144.350000 1170.500000 145.650000 ;
      RECT 1169.500000 143.650000 1186.000000 144.350000 ;
      RECT 1169.500000 142.350000 1170.500000 143.650000 ;
      RECT 0.000000 142.350000 1156.500000 145.650000 ;
      RECT 0.000000 141.650000 1170.500000 142.350000 ;
      RECT 1183.500000 140.350000 1186.000000 143.650000 ;
      RECT 1169.500000 140.350000 1170.500000 141.650000 ;
      RECT 1169.500000 139.650000 1186.000000 140.350000 ;
      RECT 1169.500000 138.350000 1170.500000 139.650000 ;
      RECT 0.000000 138.350000 1156.500000 141.650000 ;
      RECT 0.000000 137.650000 1170.500000 138.350000 ;
      RECT 1183.500000 136.350000 1186.000000 139.650000 ;
      RECT 1169.500000 136.350000 1170.500000 137.650000 ;
      RECT 1169.500000 135.650000 1186.000000 136.350000 ;
      RECT 0.000000 135.650000 1156.500000 137.650000 ;
      RECT 0.000000 135.170000 1149.500000 135.650000 ;
      RECT 1183.500000 135.165000 1186.000000 135.650000 ;
      RECT 1169.500000 134.350000 1170.500000 135.650000 ;
      RECT 1157.500000 133.650000 1170.500000 134.350000 ;
      RECT 1183.500000 132.350000 1183.980000 135.165000 ;
      RECT 1169.500000 132.350000 1170.500000 133.650000 ;
      RECT 2.020000 132.350000 1149.500000 135.170000 ;
      RECT 2.020000 132.070000 1156.500000 132.350000 ;
      RECT 1169.500000 132.065000 1183.980000 132.350000 ;
      RECT 1169.500000 131.650000 1186.000000 132.065000 ;
      RECT 1169.500000 130.350000 1170.500000 131.650000 ;
      RECT 0.000000 130.350000 1156.500000 132.070000 ;
      RECT 0.000000 129.650000 1170.500000 130.350000 ;
      RECT 1183.500000 129.485000 1186.000000 131.650000 ;
      RECT 1183.500000 128.350000 1183.980000 129.485000 ;
      RECT 1169.500000 128.350000 1170.500000 129.650000 ;
      RECT 1169.500000 127.650000 1183.980000 128.350000 ;
      RECT 1183.500000 126.385000 1183.980000 127.650000 ;
      RECT 1169.500000 126.350000 1170.500000 127.650000 ;
      RECT 0.000000 126.350000 1156.500000 129.650000 ;
      RECT 0.000000 125.650000 1170.500000 126.350000 ;
      RECT 1183.500000 125.525000 1186.000000 126.385000 ;
      RECT 0.000000 124.575000 1156.500000 125.650000 ;
      RECT 1183.500000 124.350000 1183.980000 125.525000 ;
      RECT 1169.500000 124.350000 1170.500000 125.650000 ;
      RECT 1169.500000 123.650000 1183.980000 124.350000 ;
      RECT 1183.500000 122.425000 1183.980000 123.650000 ;
      RECT 1169.500000 122.350000 1170.500000 123.650000 ;
      RECT 2.020000 122.350000 1156.500000 124.575000 ;
      RECT 2.020000 121.650000 1170.500000 122.350000 ;
      RECT 2.020000 121.475000 1156.500000 121.650000 ;
      RECT 0.000000 120.615000 1156.500000 121.475000 ;
      RECT 1183.500000 120.350000 1186.000000 122.425000 ;
      RECT 1169.500000 120.350000 1170.500000 121.650000 ;
      RECT 1169.500000 119.650000 1186.000000 120.350000 ;
      RECT 1169.500000 118.350000 1170.500000 119.650000 ;
      RECT 2.020000 118.350000 1156.500000 120.615000 ;
      RECT 2.020000 117.650000 1170.500000 118.350000 ;
      RECT 2.020000 117.515000 1156.500000 117.650000 ;
      RECT 1183.500000 116.350000 1186.000000 119.650000 ;
      RECT 1169.500000 116.350000 1170.500000 117.650000 ;
      RECT 1169.500000 115.650000 1186.000000 116.350000 ;
      RECT 0.000000 114.935000 1156.500000 117.515000 ;
      RECT 1183.500000 114.930000 1186.000000 115.650000 ;
      RECT 1169.500000 114.350000 1170.500000 115.650000 ;
      RECT 2.020000 114.350000 1156.500000 114.935000 ;
      RECT 2.020000 113.650000 1170.500000 114.350000 ;
      RECT 1183.500000 112.350000 1183.980000 114.930000 ;
      RECT 1169.500000 112.350000 1170.500000 113.650000 ;
      RECT 2.020000 111.835000 1156.500000 113.650000 ;
      RECT 1169.500000 111.830000 1183.980000 112.350000 ;
      RECT 1169.500000 111.650000 1186.000000 111.830000 ;
      RECT 1169.500000 110.350000 1170.500000 111.650000 ;
      RECT 0.000000 110.350000 1156.500000 111.835000 ;
      RECT 0.000000 109.650000 1170.500000 110.350000 ;
      RECT 1183.500000 108.350000 1186.000000 111.650000 ;
      RECT 1169.500000 108.350000 1170.500000 109.650000 ;
      RECT 1169.500000 107.650000 1186.000000 108.350000 ;
      RECT 1169.500000 106.350000 1170.500000 107.650000 ;
      RECT 0.000000 106.350000 1156.500000 109.650000 ;
      RECT 0.000000 105.650000 1170.500000 106.350000 ;
      RECT 1183.500000 104.350000 1186.000000 107.650000 ;
      RECT 1169.500000 104.350000 1170.500000 105.650000 ;
      RECT 1169.500000 103.650000 1186.000000 104.350000 ;
      RECT 1169.500000 102.350000 1170.500000 103.650000 ;
      RECT 0.000000 102.350000 1156.500000 105.650000 ;
      RECT 0.000000 101.650000 1170.500000 102.350000 ;
      RECT 1183.500000 100.350000 1186.000000 103.650000 ;
      RECT 1169.500000 100.350000 1170.500000 101.650000 ;
      RECT 1169.500000 99.650000 1186.000000 100.350000 ;
      RECT 1169.500000 98.350000 1170.500000 99.650000 ;
      RECT 0.000000 98.350000 1156.500000 101.650000 ;
      RECT 0.000000 97.650000 1170.500000 98.350000 ;
      RECT 1183.500000 96.350000 1186.000000 99.650000 ;
      RECT 1169.500000 96.350000 1170.500000 97.650000 ;
      RECT 1169.500000 95.650000 1186.000000 96.350000 ;
      RECT 1169.500000 94.350000 1170.500000 95.650000 ;
      RECT 0.000000 94.350000 1156.500000 97.650000 ;
      RECT 0.000000 93.650000 1170.500000 94.350000 ;
      RECT 1183.500000 92.350000 1186.000000 95.650000 ;
      RECT 1169.500000 92.350000 1170.500000 93.650000 ;
      RECT 1169.500000 91.650000 1186.000000 92.350000 ;
      RECT 1169.500000 90.350000 1170.500000 91.650000 ;
      RECT 0.000000 90.350000 1156.500000 93.650000 ;
      RECT 0.000000 89.650000 1170.500000 90.350000 ;
      RECT 1183.500000 88.350000 1186.000000 91.650000 ;
      RECT 1169.500000 88.350000 1170.500000 89.650000 ;
      RECT 1169.500000 87.650000 1186.000000 88.350000 ;
      RECT 1169.500000 86.350000 1170.500000 87.650000 ;
      RECT 0.000000 86.350000 1156.500000 89.650000 ;
      RECT 0.000000 85.650000 1170.500000 86.350000 ;
      RECT 1183.500000 84.350000 1186.000000 87.650000 ;
      RECT 1169.500000 84.350000 1170.500000 85.650000 ;
      RECT 1169.500000 83.650000 1186.000000 84.350000 ;
      RECT 1169.500000 82.350000 1170.500000 83.650000 ;
      RECT 0.000000 82.350000 1156.500000 85.650000 ;
      RECT 0.000000 81.650000 1170.500000 82.350000 ;
      RECT 1183.500000 80.350000 1186.000000 83.650000 ;
      RECT 1169.500000 80.350000 1170.500000 81.650000 ;
      RECT 1169.500000 79.650000 1186.000000 80.350000 ;
      RECT 1169.500000 78.350000 1170.500000 79.650000 ;
      RECT 0.000000 78.350000 1156.500000 81.650000 ;
      RECT 0.000000 77.650000 1170.500000 78.350000 ;
      RECT 1183.500000 76.350000 1186.000000 79.650000 ;
      RECT 1169.500000 76.350000 1170.500000 77.650000 ;
      RECT 1169.500000 75.650000 1186.000000 76.350000 ;
      RECT 1169.500000 74.350000 1170.500000 75.650000 ;
      RECT 0.000000 74.350000 1156.500000 77.650000 ;
      RECT 0.000000 73.650000 1170.500000 74.350000 ;
      RECT 1183.500000 72.350000 1186.000000 75.650000 ;
      RECT 1169.500000 72.350000 1170.500000 73.650000 ;
      RECT 1169.500000 71.650000 1186.000000 72.350000 ;
      RECT 1169.500000 70.350000 1170.500000 71.650000 ;
      RECT 0.000000 70.350000 1156.500000 73.650000 ;
      RECT 0.000000 69.650000 1170.500000 70.350000 ;
      RECT 1183.500000 68.350000 1186.000000 71.650000 ;
      RECT 1169.500000 68.350000 1170.500000 69.650000 ;
      RECT 1169.500000 67.650000 1186.000000 68.350000 ;
      RECT 1169.500000 66.350000 1170.500000 67.650000 ;
      RECT 0.000000 66.350000 1156.500000 69.650000 ;
      RECT 0.000000 65.650000 1170.500000 66.350000 ;
      RECT 1183.500000 64.350000 1186.000000 67.650000 ;
      RECT 1169.500000 64.350000 1170.500000 65.650000 ;
      RECT 1169.500000 63.650000 1186.000000 64.350000 ;
      RECT 1169.500000 62.350000 1170.500000 63.650000 ;
      RECT 0.000000 62.350000 1156.500000 65.650000 ;
      RECT 0.000000 61.650000 1170.500000 62.350000 ;
      RECT 1183.500000 60.350000 1186.000000 63.650000 ;
      RECT 1169.500000 60.350000 1170.500000 61.650000 ;
      RECT 1169.500000 59.650000 1186.000000 60.350000 ;
      RECT 1169.500000 58.350000 1170.500000 59.650000 ;
      RECT 0.000000 58.350000 1156.500000 61.650000 ;
      RECT 0.000000 57.650000 1170.500000 58.350000 ;
      RECT 1183.500000 56.350000 1186.000000 59.650000 ;
      RECT 1169.500000 56.350000 1170.500000 57.650000 ;
      RECT 1169.500000 55.650000 1186.000000 56.350000 ;
      RECT 1169.500000 54.350000 1170.500000 55.650000 ;
      RECT 0.000000 54.350000 1156.500000 57.650000 ;
      RECT 0.000000 53.650000 1170.500000 54.350000 ;
      RECT 1183.500000 52.350000 1186.000000 55.650000 ;
      RECT 1169.500000 52.350000 1170.500000 53.650000 ;
      RECT 1169.500000 51.650000 1186.000000 52.350000 ;
      RECT 1169.500000 50.350000 1170.500000 51.650000 ;
      RECT 0.000000 50.350000 1156.500000 53.650000 ;
      RECT 0.000000 49.650000 1170.500000 50.350000 ;
      RECT 1183.500000 48.350000 1186.000000 51.650000 ;
      RECT 1169.500000 48.350000 1170.500000 49.650000 ;
      RECT 1169.500000 47.650000 1186.000000 48.350000 ;
      RECT 0.000000 47.170000 1156.500000 49.650000 ;
      RECT 1183.500000 47.165000 1186.000000 47.650000 ;
      RECT 1169.500000 46.350000 1170.500000 47.650000 ;
      RECT 2.020000 46.350000 1156.500000 47.170000 ;
      RECT 2.020000 45.650000 1170.500000 46.350000 ;
      RECT 1183.500000 44.350000 1183.980000 47.165000 ;
      RECT 1169.500000 44.350000 1170.500000 45.650000 ;
      RECT 2.020000 44.070000 1156.500000 45.650000 ;
      RECT 1169.500000 44.065000 1183.980000 44.350000 ;
      RECT 1169.500000 43.650000 1186.000000 44.065000 ;
      RECT 1169.500000 42.350000 1170.500000 43.650000 ;
      RECT 0.000000 42.350000 1156.500000 44.070000 ;
      RECT 0.000000 41.650000 1170.500000 42.350000 ;
      RECT 1183.500000 41.485000 1186.000000 43.650000 ;
      RECT 1183.500000 40.350000 1183.980000 41.485000 ;
      RECT 1169.500000 40.350000 1170.500000 41.650000 ;
      RECT 1169.500000 39.650000 1183.980000 40.350000 ;
      RECT 1183.500000 38.385000 1183.980000 39.650000 ;
      RECT 1169.500000 38.350000 1170.500000 39.650000 ;
      RECT 0.000000 38.350000 1156.500000 41.650000 ;
      RECT 0.000000 37.650000 1170.500000 38.350000 ;
      RECT 1183.500000 37.525000 1186.000000 38.385000 ;
      RECT 0.000000 36.575000 1156.500000 37.650000 ;
      RECT 1183.500000 36.350000 1183.980000 37.525000 ;
      RECT 1169.500000 36.350000 1170.500000 37.650000 ;
      RECT 1169.500000 35.650000 1183.980000 36.350000 ;
      RECT 1183.500000 34.425000 1183.980000 35.650000 ;
      RECT 1169.500000 34.350000 1170.500000 35.650000 ;
      RECT 2.020000 34.350000 1156.500000 36.575000 ;
      RECT 2.020000 33.650000 1170.500000 34.350000 ;
      RECT 2.020000 33.475000 1156.500000 33.650000 ;
      RECT 0.000000 32.615000 1156.500000 33.475000 ;
      RECT 1183.500000 32.350000 1186.000000 34.425000 ;
      RECT 1169.500000 32.350000 1170.500000 33.650000 ;
      RECT 1169.500000 31.650000 1186.000000 32.350000 ;
      RECT 1169.500000 30.350000 1170.500000 31.650000 ;
      RECT 2.020000 30.350000 1156.500000 32.615000 ;
      RECT 2.020000 29.650000 1170.500000 30.350000 ;
      RECT 2.020000 29.515000 1156.500000 29.650000 ;
      RECT 1183.500000 28.350000 1186.000000 31.650000 ;
      RECT 1169.500000 28.350000 1170.500000 29.650000 ;
      RECT 1169.500000 27.650000 1186.000000 28.350000 ;
      RECT 0.000000 26.935000 1156.500000 29.515000 ;
      RECT 1183.500000 26.930000 1186.000000 27.650000 ;
      RECT 1169.500000 26.350000 1170.500000 27.650000 ;
      RECT 2.020000 26.350000 1156.500000 26.935000 ;
      RECT 2.020000 25.650000 1170.500000 26.350000 ;
      RECT 1183.500000 24.350000 1183.980000 26.930000 ;
      RECT 1169.500000 24.350000 1170.500000 25.650000 ;
      RECT 2.020000 23.835000 1156.500000 25.650000 ;
      RECT 1169.500000 23.830000 1183.980000 24.350000 ;
      RECT 1169.500000 23.650000 1186.000000 23.830000 ;
      RECT 1169.500000 22.350000 1170.500000 23.650000 ;
      RECT 0.000000 22.350000 1156.500000 23.835000 ;
      RECT 0.000000 21.650000 1170.500000 22.350000 ;
      RECT 1183.500000 20.350000 1186.000000 23.650000 ;
      RECT 1169.500000 20.350000 1170.500000 21.650000 ;
      RECT 1169.500000 19.650000 1186.000000 20.350000 ;
      RECT 1169.500000 18.350000 1170.500000 19.650000 ;
      RECT 0.000000 18.350000 1156.500000 21.650000 ;
      RECT 0.000000 17.650000 1170.500000 18.350000 ;
      RECT 1183.500000 16.350000 1186.000000 19.650000 ;
      RECT 1166.500000 16.350000 1170.500000 17.650000 ;
      RECT 1166.500000 15.650000 1186.000000 16.350000 ;
      RECT 1166.500000 14.350000 1170.500000 15.650000 ;
      RECT 0.000000 14.350000 1158.500000 17.650000 ;
      RECT 0.000000 13.650000 1170.500000 14.350000 ;
      RECT 1183.500000 12.350000 1186.000000 15.650000 ;
      RECT 1166.500000 12.350000 1170.500000 13.650000 ;
      RECT 1166.500000 11.650000 1186.000000 12.350000 ;
      RECT 1166.500000 10.350000 1170.500000 11.650000 ;
      RECT 0.000000 10.350000 1158.500000 13.650000 ;
      RECT 0.000000 9.650000 1170.500000 10.350000 ;
      RECT 1183.500000 8.350000 1186.000000 11.650000 ;
      RECT 1166.500000 8.350000 1170.500000 9.650000 ;
      RECT 1166.500000 7.650000 1186.000000 8.350000 ;
      RECT 1116.500000 7.650000 1158.500000 9.650000 ;
      RECT 1066.500000 7.650000 1108.500000 9.650000 ;
      RECT 1016.500000 7.650000 1058.500000 9.650000 ;
      RECT 966.500000 7.650000 1008.500000 9.650000 ;
      RECT 916.500000 7.650000 958.500000 9.650000 ;
      RECT 866.500000 7.650000 908.500000 9.650000 ;
      RECT 816.500000 7.650000 858.500000 9.650000 ;
      RECT 766.500000 7.650000 808.500000 9.650000 ;
      RECT 716.500000 7.650000 758.500000 9.650000 ;
      RECT 666.500000 7.650000 708.500000 9.650000 ;
      RECT 616.500000 7.650000 658.500000 9.650000 ;
      RECT 566.500000 7.650000 608.500000 9.650000 ;
      RECT 516.500000 7.650000 558.500000 9.650000 ;
      RECT 466.500000 7.650000 508.500000 9.650000 ;
      RECT 416.500000 7.650000 458.500000 9.650000 ;
      RECT 366.500000 7.650000 408.500000 9.650000 ;
      RECT 316.500000 7.650000 358.500000 9.650000 ;
      RECT 266.500000 7.650000 308.500000 9.650000 ;
      RECT 216.500000 7.650000 258.500000 9.650000 ;
      RECT 166.500000 7.650000 208.500000 9.650000 ;
      RECT 116.500000 7.650000 158.500000 9.650000 ;
      RECT 66.500000 7.650000 108.500000 9.650000 ;
      RECT 0.000000 7.650000 58.500000 9.650000 ;
      RECT 1166.500000 6.350000 1170.500000 7.650000 ;
      RECT 1157.500000 6.350000 1158.500000 7.650000 ;
      RECT 1116.500000 6.350000 1149.500000 7.650000 ;
      RECT 1107.500000 6.350000 1108.500000 7.650000 ;
      RECT 1066.500000 6.350000 1099.500000 7.650000 ;
      RECT 1057.500000 6.350000 1058.500000 7.650000 ;
      RECT 1016.500000 6.350000 1049.500000 7.650000 ;
      RECT 1007.500000 6.350000 1008.500000 7.650000 ;
      RECT 966.500000 6.350000 999.500000 7.650000 ;
      RECT 957.500000 6.350000 958.500000 7.650000 ;
      RECT 916.500000 6.350000 949.500000 7.650000 ;
      RECT 907.500000 6.350000 908.500000 7.650000 ;
      RECT 866.500000 6.350000 899.500000 7.650000 ;
      RECT 857.500000 6.350000 858.500000 7.650000 ;
      RECT 816.500000 6.350000 849.500000 7.650000 ;
      RECT 807.500000 6.350000 808.500000 7.650000 ;
      RECT 766.500000 6.350000 799.500000 7.650000 ;
      RECT 757.500000 6.350000 758.500000 7.650000 ;
      RECT 716.500000 6.350000 749.500000 7.650000 ;
      RECT 707.500000 6.350000 708.500000 7.650000 ;
      RECT 666.500000 6.350000 699.500000 7.650000 ;
      RECT 657.500000 6.350000 658.500000 7.650000 ;
      RECT 616.500000 6.350000 649.500000 7.650000 ;
      RECT 607.500000 6.350000 608.500000 7.650000 ;
      RECT 566.500000 6.350000 599.500000 7.650000 ;
      RECT 557.500000 6.350000 558.500000 7.650000 ;
      RECT 516.500000 6.350000 549.500000 7.650000 ;
      RECT 507.500000 6.350000 508.500000 7.650000 ;
      RECT 466.500000 6.350000 499.500000 7.650000 ;
      RECT 457.500000 6.350000 458.500000 7.650000 ;
      RECT 416.500000 6.350000 449.500000 7.650000 ;
      RECT 407.500000 6.350000 408.500000 7.650000 ;
      RECT 366.500000 6.350000 399.500000 7.650000 ;
      RECT 357.500000 6.350000 358.500000 7.650000 ;
      RECT 316.500000 6.350000 349.500000 7.650000 ;
      RECT 307.500000 6.350000 308.500000 7.650000 ;
      RECT 266.500000 6.350000 299.500000 7.650000 ;
      RECT 257.500000 6.350000 258.500000 7.650000 ;
      RECT 216.500000 6.350000 249.500000 7.650000 ;
      RECT 207.500000 6.350000 208.500000 7.650000 ;
      RECT 166.500000 6.350000 199.500000 7.650000 ;
      RECT 157.500000 6.350000 158.500000 7.650000 ;
      RECT 116.500000 6.350000 149.500000 7.650000 ;
      RECT 107.500000 6.350000 108.500000 7.650000 ;
      RECT 66.500000 6.350000 99.500000 7.650000 ;
      RECT 57.500000 6.350000 58.500000 7.650000 ;
      RECT 1157.500000 5.650000 1170.500000 6.350000 ;
      RECT 1107.500000 5.650000 1149.500000 6.350000 ;
      RECT 1057.500000 5.650000 1099.500000 6.350000 ;
      RECT 1007.500000 5.650000 1049.500000 6.350000 ;
      RECT 957.500000 5.650000 999.500000 6.350000 ;
      RECT 907.500000 5.650000 949.500000 6.350000 ;
      RECT 857.500000 5.650000 899.500000 6.350000 ;
      RECT 807.500000 5.650000 849.500000 6.350000 ;
      RECT 757.500000 5.650000 799.500000 6.350000 ;
      RECT 707.500000 5.650000 749.500000 6.350000 ;
      RECT 657.500000 5.650000 699.500000 6.350000 ;
      RECT 607.500000 5.650000 649.500000 6.350000 ;
      RECT 557.500000 5.650000 599.500000 6.350000 ;
      RECT 507.500000 5.650000 549.500000 6.350000 ;
      RECT 457.500000 5.650000 499.500000 6.350000 ;
      RECT 407.500000 5.650000 449.500000 6.350000 ;
      RECT 357.500000 5.650000 399.500000 6.350000 ;
      RECT 307.500000 5.650000 349.500000 6.350000 ;
      RECT 257.500000 5.650000 299.500000 6.350000 ;
      RECT 207.500000 5.650000 249.500000 6.350000 ;
      RECT 157.500000 5.650000 199.500000 6.350000 ;
      RECT 107.500000 5.650000 149.500000 6.350000 ;
      RECT 57.500000 5.650000 99.500000 6.350000 ;
      RECT 1183.500000 4.350000 1186.000000 7.650000 ;
      RECT 1166.500000 4.350000 1170.500000 5.650000 ;
      RECT 1157.500000 4.350000 1158.500000 5.650000 ;
      RECT 1116.500000 4.350000 1149.500000 5.650000 ;
      RECT 1107.500000 4.350000 1108.500000 5.650000 ;
      RECT 1066.500000 4.350000 1099.500000 5.650000 ;
      RECT 1057.500000 4.350000 1058.500000 5.650000 ;
      RECT 1016.500000 4.350000 1049.500000 5.650000 ;
      RECT 1007.500000 4.350000 1008.500000 5.650000 ;
      RECT 966.500000 4.350000 999.500000 5.650000 ;
      RECT 957.500000 4.350000 958.500000 5.650000 ;
      RECT 916.500000 4.350000 949.500000 5.650000 ;
      RECT 907.500000 4.350000 908.500000 5.650000 ;
      RECT 866.500000 4.350000 899.500000 5.650000 ;
      RECT 857.500000 4.350000 858.500000 5.650000 ;
      RECT 816.500000 4.350000 849.500000 5.650000 ;
      RECT 807.500000 4.350000 808.500000 5.650000 ;
      RECT 766.500000 4.350000 799.500000 5.650000 ;
      RECT 757.500000 4.350000 758.500000 5.650000 ;
      RECT 716.500000 4.350000 749.500000 5.650000 ;
      RECT 707.500000 4.350000 708.500000 5.650000 ;
      RECT 666.500000 4.350000 699.500000 5.650000 ;
      RECT 657.500000 4.350000 658.500000 5.650000 ;
      RECT 616.500000 4.350000 649.500000 5.650000 ;
      RECT 607.500000 4.350000 608.500000 5.650000 ;
      RECT 566.500000 4.350000 599.500000 5.650000 ;
      RECT 557.500000 4.350000 558.500000 5.650000 ;
      RECT 516.500000 4.350000 549.500000 5.650000 ;
      RECT 507.500000 4.350000 508.500000 5.650000 ;
      RECT 466.500000 4.350000 499.500000 5.650000 ;
      RECT 457.500000 4.350000 458.500000 5.650000 ;
      RECT 416.500000 4.350000 449.500000 5.650000 ;
      RECT 407.500000 4.350000 408.500000 5.650000 ;
      RECT 366.500000 4.350000 399.500000 5.650000 ;
      RECT 357.500000 4.350000 358.500000 5.650000 ;
      RECT 316.500000 4.350000 349.500000 5.650000 ;
      RECT 307.500000 4.350000 308.500000 5.650000 ;
      RECT 266.500000 4.350000 299.500000 5.650000 ;
      RECT 257.500000 4.350000 258.500000 5.650000 ;
      RECT 216.500000 4.350000 249.500000 5.650000 ;
      RECT 207.500000 4.350000 208.500000 5.650000 ;
      RECT 166.500000 4.350000 199.500000 5.650000 ;
      RECT 157.500000 4.350000 158.500000 5.650000 ;
      RECT 116.500000 4.350000 149.500000 5.650000 ;
      RECT 107.500000 4.350000 108.500000 5.650000 ;
      RECT 66.500000 4.350000 99.500000 5.650000 ;
      RECT 57.500000 4.350000 58.500000 5.650000 ;
      RECT 15.500000 4.350000 49.500000 7.650000 ;
      RECT 0.000000 4.350000 2.500000 7.650000 ;
      RECT 1116.500000 3.650000 1158.500000 4.350000 ;
      RECT 1066.500000 3.650000 1108.500000 4.350000 ;
      RECT 1016.500000 3.650000 1058.500000 4.350000 ;
      RECT 966.500000 3.650000 1008.500000 4.350000 ;
      RECT 916.500000 3.650000 958.500000 4.350000 ;
      RECT 866.500000 3.650000 908.500000 4.350000 ;
      RECT 816.500000 3.650000 858.500000 4.350000 ;
      RECT 766.500000 3.650000 808.500000 4.350000 ;
      RECT 716.500000 3.650000 758.500000 4.350000 ;
      RECT 666.500000 3.650000 708.500000 4.350000 ;
      RECT 616.500000 3.650000 658.500000 4.350000 ;
      RECT 566.500000 3.650000 608.500000 4.350000 ;
      RECT 516.500000 3.650000 558.500000 4.350000 ;
      RECT 466.500000 3.650000 508.500000 4.350000 ;
      RECT 416.500000 3.650000 458.500000 4.350000 ;
      RECT 366.500000 3.650000 408.500000 4.350000 ;
      RECT 316.500000 3.650000 358.500000 4.350000 ;
      RECT 266.500000 3.650000 308.500000 4.350000 ;
      RECT 216.500000 3.650000 258.500000 4.350000 ;
      RECT 166.500000 3.650000 208.500000 4.350000 ;
      RECT 116.500000 3.650000 158.500000 4.350000 ;
      RECT 66.500000 3.650000 108.500000 4.350000 ;
      RECT 0.000000 3.650000 58.500000 4.350000 ;
      RECT 1166.500000 2.350000 1186.000000 4.350000 ;
      RECT 1157.500000 2.350000 1158.500000 3.650000 ;
      RECT 1116.500000 2.350000 1149.500000 3.650000 ;
      RECT 1107.500000 2.350000 1108.500000 3.650000 ;
      RECT 1066.500000 2.350000 1099.500000 3.650000 ;
      RECT 1057.500000 2.350000 1058.500000 3.650000 ;
      RECT 1016.500000 2.350000 1049.500000 3.650000 ;
      RECT 1007.500000 2.350000 1008.500000 3.650000 ;
      RECT 966.500000 2.350000 999.500000 3.650000 ;
      RECT 957.500000 2.350000 958.500000 3.650000 ;
      RECT 916.500000 2.350000 949.500000 3.650000 ;
      RECT 907.500000 2.350000 908.500000 3.650000 ;
      RECT 866.500000 2.350000 899.500000 3.650000 ;
      RECT 857.500000 2.350000 858.500000 3.650000 ;
      RECT 816.500000 2.350000 849.500000 3.650000 ;
      RECT 807.500000 2.350000 808.500000 3.650000 ;
      RECT 766.500000 2.350000 799.500000 3.650000 ;
      RECT 757.500000 2.350000 758.500000 3.650000 ;
      RECT 716.500000 2.350000 749.500000 3.650000 ;
      RECT 707.500000 2.350000 708.500000 3.650000 ;
      RECT 666.500000 2.350000 699.500000 3.650000 ;
      RECT 657.500000 2.350000 658.500000 3.650000 ;
      RECT 616.500000 2.350000 649.500000 3.650000 ;
      RECT 607.500000 2.350000 608.500000 3.650000 ;
      RECT 566.500000 2.350000 599.500000 3.650000 ;
      RECT 557.500000 2.350000 558.500000 3.650000 ;
      RECT 516.500000 2.350000 549.500000 3.650000 ;
      RECT 507.500000 2.350000 508.500000 3.650000 ;
      RECT 466.500000 2.350000 499.500000 3.650000 ;
      RECT 457.500000 2.350000 458.500000 3.650000 ;
      RECT 416.500000 2.350000 449.500000 3.650000 ;
      RECT 407.500000 2.350000 408.500000 3.650000 ;
      RECT 366.500000 2.350000 399.500000 3.650000 ;
      RECT 357.500000 2.350000 358.500000 3.650000 ;
      RECT 316.500000 2.350000 349.500000 3.650000 ;
      RECT 307.500000 2.350000 308.500000 3.650000 ;
      RECT 266.500000 2.350000 299.500000 3.650000 ;
      RECT 257.500000 2.350000 258.500000 3.650000 ;
      RECT 216.500000 2.350000 249.500000 3.650000 ;
      RECT 207.500000 2.350000 208.500000 3.650000 ;
      RECT 166.500000 2.350000 199.500000 3.650000 ;
      RECT 157.500000 2.350000 158.500000 3.650000 ;
      RECT 116.500000 2.350000 149.500000 3.650000 ;
      RECT 107.500000 2.350000 108.500000 3.650000 ;
      RECT 66.500000 2.350000 99.500000 3.650000 ;
      RECT 57.500000 2.350000 58.500000 3.650000 ;
      RECT 857.500000 2.020000 899.500000 2.350000 ;
      RECT 807.500000 2.020000 849.500000 2.350000 ;
      RECT 757.500000 2.020000 799.500000 2.350000 ;
      RECT 707.500000 2.020000 749.500000 2.350000 ;
      RECT 607.500000 2.020000 649.500000 2.350000 ;
      RECT 557.500000 2.020000 599.500000 2.350000 ;
      RECT 507.500000 2.020000 549.500000 2.350000 ;
      RECT 457.500000 2.020000 499.500000 2.350000 ;
      RECT 357.500000 2.020000 399.500000 2.350000 ;
      RECT 257.500000 2.020000 299.500000 2.350000 ;
      RECT 107.500000 2.020000 149.500000 2.350000 ;
      RECT 1157.500000 0.350000 1186.000000 2.350000 ;
      RECT 1107.500000 0.350000 1149.500000 2.350000 ;
      RECT 1057.500000 0.350000 1099.500000 2.350000 ;
      RECT 1007.500000 0.350000 1049.500000 2.350000 ;
      RECT 957.500000 0.350000 999.500000 2.350000 ;
      RECT 907.500000 0.350000 949.500000 2.350000 ;
      RECT 899.485000 0.350000 899.500000 2.020000 ;
      RECT 857.500000 0.350000 881.830000 2.020000 ;
      RECT 819.365000 0.350000 849.500000 2.020000 ;
      RECT 799.130000 0.350000 799.500000 2.020000 ;
      RECT 757.500000 0.350000 796.030000 2.020000 ;
      RECT 733.565000 0.350000 749.500000 2.020000 ;
      RECT 707.500000 0.350000 710.230000 2.020000 ;
      RECT 657.500000 0.350000 699.500000 2.350000 ;
      RECT 647.765000 0.350000 649.500000 2.020000 ;
      RECT 607.500000 0.350000 624.430000 2.020000 ;
      RECT 561.965000 0.350000 599.500000 2.020000 ;
      RECT 557.500000 0.350000 558.865000 2.020000 ;
      RECT 507.500000 0.350000 538.630000 2.020000 ;
      RECT 476.165000 0.350000 499.500000 2.020000 ;
      RECT 457.500000 0.350000 463.425000 2.020000 ;
      RECT 407.500000 0.350000 449.500000 2.350000 ;
      RECT 390.365000 0.350000 399.500000 2.020000 ;
      RECT 357.500000 0.350000 367.030000 2.020000 ;
      RECT 307.500000 0.350000 349.500000 2.350000 ;
      RECT 298.885000 0.350000 299.500000 2.020000 ;
      RECT 257.500000 0.350000 281.230000 2.020000 ;
      RECT 207.500000 0.350000 249.500000 2.350000 ;
      RECT 157.500000 0.350000 199.500000 2.350000 ;
      RECT 132.965000 0.350000 149.500000 2.020000 ;
      RECT 107.500000 0.350000 109.630000 2.020000 ;
      RECT 57.500000 0.350000 99.500000 2.350000 ;
      RECT 0.000000 0.350000 49.500000 3.650000 ;
      RECT 905.165000 0.000000 1186.000000 0.350000 ;
      RECT 899.485000 0.000000 902.065000 0.350000 ;
      RECT 895.525000 0.000000 896.385000 2.020000 ;
      RECT 884.930000 0.000000 892.425000 2.020000 ;
      RECT 819.365000 0.000000 881.830000 0.350000 ;
      RECT 813.685000 0.000000 816.265000 2.020000 ;
      RECT 809.725000 0.000000 810.585000 2.020000 ;
      RECT 799.130000 0.000000 806.625000 0.350000 ;
      RECT 733.565000 0.000000 796.030000 0.350000 ;
      RECT 727.885000 0.000000 730.465000 2.020000 ;
      RECT 723.925000 0.000000 724.785000 2.020000 ;
      RECT 713.330000 0.000000 720.825000 2.020000 ;
      RECT 647.765000 0.000000 710.230000 0.350000 ;
      RECT 642.085000 0.000000 644.665000 2.020000 ;
      RECT 638.125000 0.000000 638.985000 2.020000 ;
      RECT 627.530000 0.000000 635.025000 2.020000 ;
      RECT 561.965000 0.000000 624.430000 0.350000 ;
      RECT 556.285000 0.000000 558.865000 0.350000 ;
      RECT 552.325000 0.000000 553.185000 0.350000 ;
      RECT 541.730000 0.000000 549.225000 2.020000 ;
      RECT 476.165000 0.000000 538.630000 0.350000 ;
      RECT 470.485000 0.000000 473.065000 2.020000 ;
      RECT 466.525000 0.000000 467.385000 2.020000 ;
      RECT 455.930000 0.000000 463.425000 0.350000 ;
      RECT 390.365000 0.000000 452.830000 0.350000 ;
      RECT 384.685000 0.000000 387.265000 2.020000 ;
      RECT 380.725000 0.000000 381.585000 2.020000 ;
      RECT 370.130000 0.000000 377.625000 2.020000 ;
      RECT 304.565000 0.000000 367.030000 0.350000 ;
      RECT 298.885000 0.000000 301.465000 0.350000 ;
      RECT 294.925000 0.000000 295.785000 2.020000 ;
      RECT 284.330000 0.000000 291.825000 2.020000 ;
      RECT 132.965000 0.000000 281.230000 0.350000 ;
      RECT 127.285000 0.000000 129.865000 2.020000 ;
      RECT 123.325000 0.000000 124.185000 2.020000 ;
      RECT 112.730000 0.000000 120.225000 2.020000 ;
      RECT 0.000000 0.000000 109.630000 0.350000 ;
    LAYER M3 ;
      RECT 1139.000000 685.650000 1186.000000 686.000000 ;
      RECT 0.000000 685.650000 670.000000 686.000000 ;
      RECT 1139.000000 683.650000 1158.500000 685.650000 ;
      RECT 616.500000 683.650000 658.500000 685.650000 ;
      RECT 566.500000 683.650000 608.500000 685.650000 ;
      RECT 516.500000 683.650000 558.500000 685.650000 ;
      RECT 466.500000 683.650000 508.500000 685.650000 ;
      RECT 416.500000 683.650000 458.500000 685.650000 ;
      RECT 366.500000 683.650000 408.500000 685.650000 ;
      RECT 316.500000 683.650000 358.500000 685.650000 ;
      RECT 0.000000 683.650000 308.500000 685.650000 ;
      RECT 1166.500000 682.350000 1186.000000 685.650000 ;
      RECT 1157.500000 682.350000 1158.500000 683.650000 ;
      RECT 666.500000 682.350000 670.000000 685.650000 ;
      RECT 657.500000 682.350000 658.500000 683.650000 ;
      RECT 616.500000 682.350000 649.500000 683.650000 ;
      RECT 607.500000 682.350000 608.500000 683.650000 ;
      RECT 566.500000 682.350000 599.500000 683.650000 ;
      RECT 557.500000 682.350000 558.500000 683.650000 ;
      RECT 516.500000 682.350000 549.500000 683.650000 ;
      RECT 507.500000 682.350000 508.500000 683.650000 ;
      RECT 466.500000 682.350000 499.500000 683.650000 ;
      RECT 457.500000 682.350000 458.500000 683.650000 ;
      RECT 416.500000 682.350000 449.500000 683.650000 ;
      RECT 407.500000 682.350000 408.500000 683.650000 ;
      RECT 366.500000 682.350000 383.500000 683.650000 ;
      RECT 357.500000 682.350000 358.500000 683.650000 ;
      RECT 316.500000 682.350000 349.500000 683.650000 ;
      RECT 307.500000 682.350000 308.500000 683.650000 ;
      RECT 1157.500000 681.650000 1186.000000 682.350000 ;
      RECT 657.500000 681.650000 670.000000 682.350000 ;
      RECT 607.500000 681.650000 649.500000 682.350000 ;
      RECT 557.500000 681.650000 599.500000 682.350000 ;
      RECT 507.500000 681.650000 549.500000 682.350000 ;
      RECT 457.500000 681.650000 499.500000 682.350000 ;
      RECT 407.500000 681.650000 449.500000 682.350000 ;
      RECT 357.500000 681.650000 383.500000 682.350000 ;
      RECT 307.500000 681.650000 349.500000 682.350000 ;
      RECT 1157.500000 680.350000 1158.500000 681.650000 ;
      RECT 1139.000000 680.350000 1149.500000 683.650000 ;
      RECT 657.500000 680.350000 658.500000 681.650000 ;
      RECT 616.500000 680.350000 649.500000 681.650000 ;
      RECT 607.500000 680.350000 608.500000 681.650000 ;
      RECT 566.500000 680.350000 599.500000 681.650000 ;
      RECT 557.500000 680.350000 558.500000 681.650000 ;
      RECT 516.500000 680.350000 549.500000 681.650000 ;
      RECT 507.500000 680.350000 508.500000 681.650000 ;
      RECT 466.500000 680.350000 499.500000 681.650000 ;
      RECT 457.500000 680.350000 458.500000 681.650000 ;
      RECT 416.500000 680.350000 449.500000 681.650000 ;
      RECT 407.500000 680.350000 408.500000 681.650000 ;
      RECT 396.500000 680.350000 399.500000 683.650000 ;
      RECT 366.500000 680.350000 383.500000 681.650000 ;
      RECT 357.500000 680.350000 358.500000 681.650000 ;
      RECT 316.500000 680.350000 349.500000 681.650000 ;
      RECT 307.500000 680.350000 308.500000 681.650000 ;
      RECT 0.000000 680.350000 299.500000 683.650000 ;
      RECT 1139.000000 679.650000 1158.500000 680.350000 ;
      RECT 616.500000 679.650000 658.500000 680.350000 ;
      RECT 566.500000 679.650000 608.500000 680.350000 ;
      RECT 516.500000 679.650000 558.500000 680.350000 ;
      RECT 466.500000 679.650000 508.500000 680.350000 ;
      RECT 416.500000 679.650000 458.500000 680.350000 ;
      RECT 366.500000 679.650000 408.500000 680.350000 ;
      RECT 316.500000 679.650000 358.500000 680.350000 ;
      RECT 0.000000 679.650000 308.500000 680.350000 ;
      RECT 1166.500000 678.350000 1186.000000 681.650000 ;
      RECT 1157.500000 678.350000 1158.500000 679.650000 ;
      RECT 666.500000 678.350000 670.000000 681.650000 ;
      RECT 657.500000 678.350000 658.500000 679.650000 ;
      RECT 616.500000 678.350000 649.500000 679.650000 ;
      RECT 607.500000 678.350000 608.500000 679.650000 ;
      RECT 566.500000 678.350000 599.500000 679.650000 ;
      RECT 557.500000 678.350000 558.500000 679.650000 ;
      RECT 516.500000 678.350000 549.500000 679.650000 ;
      RECT 507.500000 678.350000 508.500000 679.650000 ;
      RECT 466.500000 678.350000 499.500000 679.650000 ;
      RECT 457.500000 678.350000 458.500000 679.650000 ;
      RECT 416.500000 678.350000 449.500000 679.650000 ;
      RECT 407.500000 678.350000 408.500000 679.650000 ;
      RECT 366.500000 678.350000 383.500000 679.650000 ;
      RECT 357.500000 678.350000 358.500000 679.650000 ;
      RECT 316.500000 678.350000 349.500000 679.650000 ;
      RECT 307.500000 678.350000 308.500000 679.650000 ;
      RECT 1157.500000 677.650000 1186.000000 678.350000 ;
      RECT 657.500000 677.650000 670.000000 678.350000 ;
      RECT 607.500000 677.650000 649.500000 678.350000 ;
      RECT 557.500000 677.650000 599.500000 678.350000 ;
      RECT 507.500000 677.650000 549.500000 678.350000 ;
      RECT 457.500000 677.650000 499.500000 678.350000 ;
      RECT 407.500000 677.650000 449.500000 678.350000 ;
      RECT 357.500000 677.650000 383.500000 678.350000 ;
      RECT 1157.500000 676.350000 1158.500000 677.650000 ;
      RECT 1139.000000 676.350000 1149.500000 679.650000 ;
      RECT 657.500000 676.350000 658.500000 677.650000 ;
      RECT 616.500000 676.350000 649.500000 677.650000 ;
      RECT 607.500000 676.350000 608.500000 677.650000 ;
      RECT 566.500000 676.350000 599.500000 677.650000 ;
      RECT 557.500000 676.350000 558.500000 677.650000 ;
      RECT 516.500000 676.350000 549.500000 677.650000 ;
      RECT 507.500000 676.350000 508.500000 677.650000 ;
      RECT 466.500000 676.350000 499.500000 677.650000 ;
      RECT 457.500000 676.350000 458.500000 677.650000 ;
      RECT 416.500000 676.350000 449.500000 677.650000 ;
      RECT 407.500000 676.350000 408.500000 677.650000 ;
      RECT 396.500000 676.350000 399.500000 679.650000 ;
      RECT 366.500000 676.350000 383.500000 677.650000 ;
      RECT 357.500000 676.350000 358.500000 677.650000 ;
      RECT 307.500000 676.350000 349.500000 678.350000 ;
      RECT 0.000000 676.350000 299.500000 679.650000 ;
      RECT 1139.000000 675.650000 1158.500000 676.350000 ;
      RECT 616.500000 675.650000 658.500000 676.350000 ;
      RECT 566.500000 675.650000 608.500000 676.350000 ;
      RECT 516.500000 675.650000 558.500000 676.350000 ;
      RECT 466.500000 675.650000 508.500000 676.350000 ;
      RECT 416.500000 675.650000 458.500000 676.350000 ;
      RECT 366.500000 675.650000 408.500000 676.350000 ;
      RECT 0.000000 675.650000 358.500000 676.350000 ;
      RECT 1166.500000 674.350000 1186.000000 677.650000 ;
      RECT 1157.500000 674.350000 1158.500000 675.650000 ;
      RECT 666.500000 674.350000 670.000000 677.650000 ;
      RECT 657.500000 674.350000 658.500000 675.650000 ;
      RECT 616.500000 674.350000 649.500000 675.650000 ;
      RECT 607.500000 674.350000 608.500000 675.650000 ;
      RECT 566.500000 674.350000 599.500000 675.650000 ;
      RECT 557.500000 674.350000 558.500000 675.650000 ;
      RECT 516.500000 674.350000 549.500000 675.650000 ;
      RECT 507.500000 674.350000 508.500000 675.650000 ;
      RECT 466.500000 674.350000 499.500000 675.650000 ;
      RECT 457.500000 674.350000 458.500000 675.650000 ;
      RECT 416.500000 674.350000 449.500000 675.650000 ;
      RECT 407.500000 674.350000 408.500000 675.650000 ;
      RECT 366.500000 674.350000 383.500000 675.650000 ;
      RECT 357.500000 674.350000 358.500000 675.650000 ;
      RECT 1157.500000 673.650000 1186.000000 674.350000 ;
      RECT 657.500000 673.650000 670.000000 674.350000 ;
      RECT 607.500000 673.650000 649.500000 674.350000 ;
      RECT 557.500000 673.650000 599.500000 674.350000 ;
      RECT 507.500000 673.650000 549.500000 674.350000 ;
      RECT 457.500000 673.650000 499.500000 674.350000 ;
      RECT 407.500000 673.650000 449.500000 674.350000 ;
      RECT 357.500000 673.650000 383.500000 674.350000 ;
      RECT 1157.500000 672.350000 1158.500000 673.650000 ;
      RECT 1139.000000 672.350000 1149.500000 675.650000 ;
      RECT 657.500000 672.350000 658.500000 673.650000 ;
      RECT 616.500000 672.350000 649.500000 673.650000 ;
      RECT 607.500000 672.350000 608.500000 673.650000 ;
      RECT 566.500000 672.350000 599.500000 673.650000 ;
      RECT 557.500000 672.350000 558.500000 673.650000 ;
      RECT 516.500000 672.350000 549.500000 673.650000 ;
      RECT 507.500000 672.350000 508.500000 673.650000 ;
      RECT 466.500000 672.350000 499.500000 673.650000 ;
      RECT 457.500000 672.350000 458.500000 673.650000 ;
      RECT 416.500000 672.350000 449.500000 673.650000 ;
      RECT 407.500000 672.350000 408.500000 673.650000 ;
      RECT 396.500000 672.350000 399.500000 675.650000 ;
      RECT 366.500000 672.350000 383.500000 673.650000 ;
      RECT 357.500000 672.350000 358.500000 673.650000 ;
      RECT 0.000000 672.350000 349.500000 675.650000 ;
      RECT 1139.000000 671.650000 1158.500000 672.350000 ;
      RECT 616.500000 671.650000 658.500000 672.350000 ;
      RECT 566.500000 671.650000 608.500000 672.350000 ;
      RECT 516.500000 671.650000 558.500000 672.350000 ;
      RECT 466.500000 671.650000 508.500000 672.350000 ;
      RECT 416.500000 671.650000 458.500000 672.350000 ;
      RECT 366.500000 671.650000 408.500000 672.350000 ;
      RECT 0.000000 671.650000 358.500000 672.350000 ;
      RECT 1166.500000 670.350000 1186.000000 673.650000 ;
      RECT 1157.500000 670.350000 1158.500000 671.650000 ;
      RECT 666.500000 670.350000 670.000000 673.650000 ;
      RECT 657.500000 670.350000 658.500000 671.650000 ;
      RECT 616.500000 670.350000 649.500000 671.650000 ;
      RECT 607.500000 670.350000 608.500000 671.650000 ;
      RECT 566.500000 670.350000 599.500000 671.650000 ;
      RECT 557.500000 670.350000 558.500000 671.650000 ;
      RECT 516.500000 670.350000 549.500000 671.650000 ;
      RECT 507.500000 670.350000 508.500000 671.650000 ;
      RECT 466.500000 670.350000 499.500000 671.650000 ;
      RECT 457.500000 670.350000 458.500000 671.650000 ;
      RECT 416.500000 670.350000 449.500000 671.650000 ;
      RECT 407.500000 670.350000 408.500000 671.650000 ;
      RECT 366.500000 670.350000 383.500000 671.650000 ;
      RECT 357.500000 670.350000 358.500000 671.650000 ;
      RECT 1157.500000 669.650000 1186.000000 670.350000 ;
      RECT 657.500000 669.650000 670.000000 670.350000 ;
      RECT 607.500000 669.650000 649.500000 670.350000 ;
      RECT 557.500000 669.650000 599.500000 670.350000 ;
      RECT 507.500000 669.650000 549.500000 670.350000 ;
      RECT 457.500000 669.650000 499.500000 670.350000 ;
      RECT 407.500000 669.650000 449.500000 670.350000 ;
      RECT 357.500000 669.650000 383.500000 670.350000 ;
      RECT 1157.500000 668.350000 1158.500000 669.650000 ;
      RECT 1139.000000 668.350000 1149.500000 671.650000 ;
      RECT 657.500000 668.350000 658.500000 669.650000 ;
      RECT 616.500000 668.350000 649.500000 669.650000 ;
      RECT 607.500000 668.350000 608.500000 669.650000 ;
      RECT 566.500000 668.350000 599.500000 669.650000 ;
      RECT 557.500000 668.350000 558.500000 669.650000 ;
      RECT 516.500000 668.350000 549.500000 669.650000 ;
      RECT 507.500000 668.350000 508.500000 669.650000 ;
      RECT 466.500000 668.350000 499.500000 669.650000 ;
      RECT 457.500000 668.350000 458.500000 669.650000 ;
      RECT 416.500000 668.350000 449.500000 669.650000 ;
      RECT 407.500000 668.350000 408.500000 669.650000 ;
      RECT 396.500000 668.350000 399.500000 671.650000 ;
      RECT 382.500000 668.350000 383.500000 669.650000 ;
      RECT 357.500000 668.350000 358.500000 669.650000 ;
      RECT 0.000000 668.350000 349.500000 671.650000 ;
      RECT 1139.000000 667.650000 1158.500000 668.350000 ;
      RECT 616.500000 667.650000 658.500000 668.350000 ;
      RECT 566.500000 667.650000 608.500000 668.350000 ;
      RECT 516.500000 667.650000 558.500000 668.350000 ;
      RECT 466.500000 667.650000 508.500000 668.350000 ;
      RECT 416.500000 667.650000 458.500000 668.350000 ;
      RECT 382.500000 667.650000 408.500000 668.350000 ;
      RECT 0.000000 667.650000 358.500000 668.350000 ;
      RECT 1166.500000 666.350000 1186.000000 669.650000 ;
      RECT 1157.500000 666.350000 1158.500000 667.650000 ;
      RECT 666.500000 666.350000 670.000000 669.650000 ;
      RECT 657.500000 666.350000 658.500000 667.650000 ;
      RECT 616.500000 666.350000 649.500000 667.650000 ;
      RECT 607.500000 666.350000 608.500000 667.650000 ;
      RECT 566.500000 666.350000 599.500000 667.650000 ;
      RECT 557.500000 666.350000 558.500000 667.650000 ;
      RECT 516.500000 666.350000 549.500000 667.650000 ;
      RECT 507.500000 666.350000 508.500000 667.650000 ;
      RECT 466.500000 666.350000 499.500000 667.650000 ;
      RECT 457.500000 666.350000 458.500000 667.650000 ;
      RECT 416.500000 666.350000 449.500000 667.650000 ;
      RECT 407.500000 666.350000 408.500000 667.650000 ;
      RECT 382.500000 666.350000 383.500000 667.650000 ;
      RECT 366.500000 666.350000 369.500000 669.650000 ;
      RECT 357.500000 666.350000 358.500000 667.650000 ;
      RECT 1157.500000 665.650000 1186.000000 666.350000 ;
      RECT 657.500000 665.650000 670.000000 666.350000 ;
      RECT 607.500000 665.650000 649.500000 666.350000 ;
      RECT 557.500000 665.650000 599.500000 666.350000 ;
      RECT 507.500000 665.650000 549.500000 666.350000 ;
      RECT 457.500000 665.650000 499.500000 666.350000 ;
      RECT 407.500000 665.650000 449.500000 666.350000 ;
      RECT 357.500000 665.650000 383.500000 666.350000 ;
      RECT 1157.500000 664.350000 1158.500000 665.650000 ;
      RECT 1139.000000 664.350000 1149.500000 667.650000 ;
      RECT 657.500000 664.350000 658.500000 665.650000 ;
      RECT 616.500000 664.350000 649.500000 665.650000 ;
      RECT 607.500000 664.350000 608.500000 665.650000 ;
      RECT 566.500000 664.350000 599.500000 665.650000 ;
      RECT 557.500000 664.350000 558.500000 665.650000 ;
      RECT 516.500000 664.350000 549.500000 665.650000 ;
      RECT 507.500000 664.350000 508.500000 665.650000 ;
      RECT 466.500000 664.350000 499.500000 665.650000 ;
      RECT 457.500000 664.350000 458.500000 665.650000 ;
      RECT 416.500000 664.350000 449.500000 665.650000 ;
      RECT 407.500000 664.350000 408.500000 665.650000 ;
      RECT 396.500000 664.350000 399.500000 667.650000 ;
      RECT 382.500000 664.350000 383.500000 665.650000 ;
      RECT 357.500000 664.350000 358.500000 665.650000 ;
      RECT 0.000000 664.350000 349.500000 667.650000 ;
      RECT 1139.000000 663.650000 1158.500000 664.350000 ;
      RECT 616.500000 663.650000 658.500000 664.350000 ;
      RECT 566.500000 663.650000 608.500000 664.350000 ;
      RECT 516.500000 663.650000 558.500000 664.350000 ;
      RECT 466.500000 663.650000 508.500000 664.350000 ;
      RECT 416.500000 663.650000 458.500000 664.350000 ;
      RECT 382.500000 663.650000 408.500000 664.350000 ;
      RECT 0.000000 663.650000 358.500000 664.350000 ;
      RECT 1166.500000 662.350000 1186.000000 665.650000 ;
      RECT 1157.500000 662.350000 1158.500000 663.650000 ;
      RECT 666.500000 662.350000 670.000000 665.650000 ;
      RECT 657.500000 662.350000 658.500000 663.650000 ;
      RECT 616.500000 662.350000 649.500000 663.650000 ;
      RECT 607.500000 662.350000 608.500000 663.650000 ;
      RECT 566.500000 662.350000 599.500000 663.650000 ;
      RECT 557.500000 662.350000 558.500000 663.650000 ;
      RECT 516.500000 662.350000 549.500000 663.650000 ;
      RECT 507.500000 662.350000 508.500000 663.650000 ;
      RECT 466.500000 662.350000 499.500000 663.650000 ;
      RECT 457.500000 662.350000 458.500000 663.650000 ;
      RECT 416.500000 662.350000 449.500000 663.650000 ;
      RECT 407.500000 662.350000 408.500000 663.650000 ;
      RECT 382.500000 662.350000 383.500000 663.650000 ;
      RECT 366.500000 662.350000 369.500000 665.650000 ;
      RECT 357.500000 662.350000 358.500000 663.650000 ;
      RECT 1157.500000 661.650000 1186.000000 662.350000 ;
      RECT 657.500000 661.650000 670.000000 662.350000 ;
      RECT 607.500000 661.650000 649.500000 662.350000 ;
      RECT 557.500000 661.650000 599.500000 662.350000 ;
      RECT 507.500000 661.650000 549.500000 662.350000 ;
      RECT 457.500000 661.650000 499.500000 662.350000 ;
      RECT 407.500000 661.650000 449.500000 662.350000 ;
      RECT 357.500000 661.650000 383.500000 662.350000 ;
      RECT 1157.500000 660.350000 1158.500000 661.650000 ;
      RECT 1139.000000 660.350000 1149.500000 663.650000 ;
      RECT 657.500000 660.350000 658.500000 661.650000 ;
      RECT 616.500000 660.350000 649.500000 661.650000 ;
      RECT 607.500000 660.350000 608.500000 661.650000 ;
      RECT 566.500000 660.350000 599.500000 661.650000 ;
      RECT 557.500000 660.350000 558.500000 661.650000 ;
      RECT 516.500000 660.350000 549.500000 661.650000 ;
      RECT 507.500000 660.350000 508.500000 661.650000 ;
      RECT 466.500000 660.350000 499.500000 661.650000 ;
      RECT 457.500000 660.350000 458.500000 661.650000 ;
      RECT 416.500000 660.350000 449.500000 661.650000 ;
      RECT 407.500000 660.350000 408.500000 661.650000 ;
      RECT 396.500000 660.350000 399.500000 663.650000 ;
      RECT 382.500000 660.350000 383.500000 661.650000 ;
      RECT 357.500000 660.350000 358.500000 661.650000 ;
      RECT 0.000000 660.350000 349.500000 663.650000 ;
      RECT 1139.000000 659.650000 1158.500000 660.350000 ;
      RECT 616.500000 659.650000 658.500000 660.350000 ;
      RECT 566.500000 659.650000 608.500000 660.350000 ;
      RECT 516.500000 659.650000 558.500000 660.350000 ;
      RECT 466.500000 659.650000 508.500000 660.350000 ;
      RECT 416.500000 659.650000 458.500000 660.350000 ;
      RECT 382.500000 659.650000 408.500000 660.350000 ;
      RECT 0.000000 659.650000 358.500000 660.350000 ;
      RECT 1166.500000 658.350000 1186.000000 661.650000 ;
      RECT 1157.500000 658.350000 1158.500000 659.650000 ;
      RECT 666.500000 658.350000 670.000000 661.650000 ;
      RECT 657.500000 658.350000 658.500000 659.650000 ;
      RECT 616.500000 658.350000 649.500000 659.650000 ;
      RECT 607.500000 658.350000 608.500000 659.650000 ;
      RECT 566.500000 658.350000 599.500000 659.650000 ;
      RECT 557.500000 658.350000 558.500000 659.650000 ;
      RECT 516.500000 658.350000 549.500000 659.650000 ;
      RECT 507.500000 658.350000 508.500000 659.650000 ;
      RECT 466.500000 658.350000 499.500000 659.650000 ;
      RECT 457.500000 658.350000 458.500000 659.650000 ;
      RECT 416.500000 658.350000 449.500000 659.650000 ;
      RECT 407.500000 658.350000 408.500000 659.650000 ;
      RECT 382.500000 658.350000 383.500000 659.650000 ;
      RECT 366.500000 658.350000 369.500000 661.650000 ;
      RECT 357.500000 658.350000 358.500000 659.650000 ;
      RECT 1157.500000 657.650000 1186.000000 658.350000 ;
      RECT 357.500000 657.650000 383.500000 658.350000 ;
      RECT 1157.500000 656.350000 1158.500000 657.650000 ;
      RECT 1139.000000 656.350000 1149.500000 659.650000 ;
      RECT 657.500000 656.350000 670.000000 658.350000 ;
      RECT 607.500000 656.350000 649.500000 658.350000 ;
      RECT 557.500000 656.350000 599.500000 658.350000 ;
      RECT 507.500000 656.350000 549.500000 658.350000 ;
      RECT 457.500000 656.350000 499.500000 658.350000 ;
      RECT 407.500000 656.350000 449.500000 658.350000 ;
      RECT 396.500000 656.350000 399.500000 659.650000 ;
      RECT 382.500000 656.350000 383.500000 657.650000 ;
      RECT 357.500000 656.350000 358.500000 657.650000 ;
      RECT 0.000000 656.350000 349.500000 659.650000 ;
      RECT 382.500000 656.000000 670.000000 656.350000 ;
      RECT 1139.000000 655.650000 1158.500000 656.350000 ;
      RECT 382.500000 655.650000 399.000000 656.000000 ;
      RECT 0.000000 655.650000 358.500000 656.350000 ;
      RECT 1166.500000 654.350000 1186.000000 657.650000 ;
      RECT 1157.500000 654.350000 1158.500000 655.650000 ;
      RECT 382.500000 654.350000 383.500000 655.650000 ;
      RECT 366.500000 654.350000 369.500000 657.650000 ;
      RECT 357.500000 654.350000 358.500000 655.650000 ;
      RECT 1157.500000 653.650000 1186.000000 654.350000 ;
      RECT 357.500000 653.650000 383.500000 654.350000 ;
      RECT 1157.500000 652.350000 1158.500000 653.650000 ;
      RECT 1139.000000 652.350000 1149.500000 655.650000 ;
      RECT 396.500000 652.350000 399.000000 655.650000 ;
      RECT 382.500000 652.350000 383.500000 653.650000 ;
      RECT 357.500000 652.350000 358.500000 653.650000 ;
      RECT 0.000000 652.350000 349.500000 655.650000 ;
      RECT 1139.000000 651.650000 1158.500000 652.350000 ;
      RECT 382.500000 651.650000 399.000000 652.350000 ;
      RECT 0.000000 651.650000 358.500000 652.350000 ;
      RECT 1166.500000 650.350000 1186.000000 653.650000 ;
      RECT 1157.500000 650.350000 1158.500000 651.650000 ;
      RECT 382.500000 650.350000 383.500000 651.650000 ;
      RECT 366.500000 650.350000 369.500000 653.650000 ;
      RECT 357.500000 650.350000 358.500000 651.650000 ;
      RECT 1157.500000 649.650000 1186.000000 650.350000 ;
      RECT 357.500000 649.650000 383.500000 650.350000 ;
      RECT 1157.500000 648.350000 1158.500000 649.650000 ;
      RECT 1139.000000 648.350000 1149.500000 651.650000 ;
      RECT 396.500000 648.350000 399.000000 651.650000 ;
      RECT 382.500000 648.350000 383.500000 649.650000 ;
      RECT 357.500000 648.350000 358.500000 649.650000 ;
      RECT 0.000000 648.350000 349.500000 651.650000 ;
      RECT 1139.000000 647.650000 1158.500000 648.350000 ;
      RECT 382.500000 647.650000 399.000000 648.350000 ;
      RECT 0.000000 647.650000 358.500000 648.350000 ;
      RECT 1166.500000 646.350000 1186.000000 649.650000 ;
      RECT 1157.500000 646.350000 1158.500000 647.650000 ;
      RECT 382.500000 646.350000 383.500000 647.650000 ;
      RECT 366.500000 646.350000 369.500000 649.650000 ;
      RECT 357.500000 646.350000 358.500000 647.650000 ;
      RECT 1157.500000 645.650000 1186.000000 646.350000 ;
      RECT 357.500000 645.650000 383.500000 646.350000 ;
      RECT 1157.500000 644.350000 1158.500000 645.650000 ;
      RECT 1139.000000 644.350000 1149.500000 647.650000 ;
      RECT 396.500000 644.350000 399.000000 647.650000 ;
      RECT 382.500000 644.350000 383.500000 645.650000 ;
      RECT 357.500000 644.350000 358.500000 645.650000 ;
      RECT 0.000000 644.350000 349.500000 647.650000 ;
      RECT 1139.000000 643.650000 1158.500000 644.350000 ;
      RECT 382.500000 643.650000 399.000000 644.350000 ;
      RECT 0.000000 643.650000 358.500000 644.350000 ;
      RECT 1166.500000 642.350000 1186.000000 645.650000 ;
      RECT 1157.500000 642.350000 1158.500000 643.650000 ;
      RECT 382.500000 642.350000 383.500000 643.650000 ;
      RECT 366.500000 642.350000 369.500000 645.650000 ;
      RECT 357.500000 642.350000 358.500000 643.650000 ;
      RECT 1157.500000 641.650000 1186.000000 642.350000 ;
      RECT 357.500000 641.650000 383.500000 642.350000 ;
      RECT 1157.500000 640.350000 1158.500000 641.650000 ;
      RECT 1139.000000 640.350000 1149.500000 643.650000 ;
      RECT 396.500000 640.350000 399.000000 643.650000 ;
      RECT 382.500000 640.350000 383.500000 641.650000 ;
      RECT 357.500000 640.350000 358.500000 641.650000 ;
      RECT 0.000000 640.350000 349.500000 643.650000 ;
      RECT 1139.000000 639.650000 1158.500000 640.350000 ;
      RECT 382.500000 639.650000 399.000000 640.350000 ;
      RECT 0.000000 639.650000 358.500000 640.350000 ;
      RECT 1166.500000 638.350000 1186.000000 641.650000 ;
      RECT 1157.500000 638.350000 1158.500000 639.650000 ;
      RECT 382.500000 638.350000 383.500000 639.650000 ;
      RECT 366.500000 638.350000 369.500000 641.650000 ;
      RECT 357.500000 638.350000 358.500000 639.650000 ;
      RECT 1157.500000 637.650000 1186.000000 638.350000 ;
      RECT 357.500000 637.650000 383.500000 638.350000 ;
      RECT 1157.500000 636.350000 1158.500000 637.650000 ;
      RECT 1139.000000 636.350000 1149.500000 639.650000 ;
      RECT 396.500000 636.350000 399.000000 639.650000 ;
      RECT 382.500000 636.350000 383.500000 637.650000 ;
      RECT 357.500000 636.350000 358.500000 637.650000 ;
      RECT 0.000000 636.350000 349.500000 639.650000 ;
      RECT 1139.000000 635.650000 1158.500000 636.350000 ;
      RECT 382.500000 635.650000 399.000000 636.350000 ;
      RECT 0.000000 635.650000 358.500000 636.350000 ;
      RECT 1166.500000 634.350000 1186.000000 637.650000 ;
      RECT 1157.500000 634.350000 1158.500000 635.650000 ;
      RECT 382.500000 634.350000 383.500000 635.650000 ;
      RECT 366.500000 634.350000 369.500000 637.650000 ;
      RECT 357.500000 634.350000 358.500000 635.650000 ;
      RECT 1157.500000 633.650000 1186.000000 634.350000 ;
      RECT 357.500000 633.650000 383.500000 634.350000 ;
      RECT 1157.500000 632.350000 1158.500000 633.650000 ;
      RECT 1139.000000 632.350000 1149.500000 635.650000 ;
      RECT 396.500000 632.350000 399.000000 635.650000 ;
      RECT 382.500000 632.350000 383.500000 633.650000 ;
      RECT 357.500000 632.350000 358.500000 633.650000 ;
      RECT 0.000000 632.350000 349.500000 635.650000 ;
      RECT 1139.000000 631.650000 1158.500000 632.350000 ;
      RECT 382.500000 631.650000 399.000000 632.350000 ;
      RECT 0.000000 631.650000 358.500000 632.350000 ;
      RECT 1166.500000 630.350000 1186.000000 633.650000 ;
      RECT 1157.500000 630.350000 1158.500000 631.650000 ;
      RECT 382.500000 630.350000 383.500000 631.650000 ;
      RECT 366.500000 630.350000 369.500000 633.650000 ;
      RECT 357.500000 630.350000 358.500000 631.650000 ;
      RECT 1157.500000 629.650000 1186.000000 630.350000 ;
      RECT 357.500000 629.650000 383.500000 630.350000 ;
      RECT 1157.500000 628.350000 1158.500000 629.650000 ;
      RECT 1139.000000 628.350000 1149.500000 631.650000 ;
      RECT 396.500000 628.350000 399.000000 631.650000 ;
      RECT 382.500000 628.350000 383.500000 629.650000 ;
      RECT 357.500000 628.350000 358.500000 629.650000 ;
      RECT 0.000000 628.350000 349.500000 631.650000 ;
      RECT 1139.000000 627.650000 1158.500000 628.350000 ;
      RECT 382.500000 627.650000 399.000000 628.350000 ;
      RECT 0.000000 627.650000 358.500000 628.350000 ;
      RECT 1166.500000 626.350000 1186.000000 629.650000 ;
      RECT 1157.500000 626.350000 1158.500000 627.650000 ;
      RECT 382.500000 626.350000 383.500000 627.650000 ;
      RECT 366.500000 626.350000 369.500000 629.650000 ;
      RECT 357.500000 626.350000 358.500000 627.650000 ;
      RECT 1157.500000 625.650000 1186.000000 626.350000 ;
      RECT 357.500000 625.650000 383.500000 626.350000 ;
      RECT 1157.500000 624.350000 1158.500000 625.650000 ;
      RECT 1139.000000 624.350000 1149.500000 627.650000 ;
      RECT 396.500000 624.350000 399.000000 627.650000 ;
      RECT 382.500000 624.350000 383.500000 625.650000 ;
      RECT 357.500000 624.350000 358.500000 625.650000 ;
      RECT 0.000000 624.350000 349.500000 627.650000 ;
      RECT 1139.000000 623.650000 1158.500000 624.350000 ;
      RECT 382.500000 623.650000 399.000000 624.350000 ;
      RECT 0.000000 623.650000 358.500000 624.350000 ;
      RECT 1166.500000 622.350000 1186.000000 625.650000 ;
      RECT 1157.500000 622.350000 1158.500000 623.650000 ;
      RECT 382.500000 622.350000 383.500000 623.650000 ;
      RECT 366.500000 622.350000 369.500000 625.650000 ;
      RECT 357.500000 622.350000 358.500000 623.650000 ;
      RECT 1157.500000 621.650000 1186.000000 622.350000 ;
      RECT 357.500000 621.650000 383.500000 622.350000 ;
      RECT 1157.500000 620.350000 1158.500000 621.650000 ;
      RECT 1139.000000 620.350000 1149.500000 623.650000 ;
      RECT 396.500000 620.350000 399.000000 623.650000 ;
      RECT 382.500000 620.350000 383.500000 621.650000 ;
      RECT 357.500000 620.350000 358.500000 621.650000 ;
      RECT 0.000000 620.350000 349.500000 623.650000 ;
      RECT 1139.000000 619.650000 1158.500000 620.350000 ;
      RECT 382.500000 619.650000 399.000000 620.350000 ;
      RECT 0.000000 619.650000 358.500000 620.350000 ;
      RECT 1166.500000 618.350000 1186.000000 621.650000 ;
      RECT 1157.500000 618.350000 1158.500000 619.650000 ;
      RECT 382.500000 618.350000 383.500000 619.650000 ;
      RECT 366.500000 618.350000 369.500000 621.650000 ;
      RECT 357.500000 618.350000 358.500000 619.650000 ;
      RECT 1157.500000 617.650000 1186.000000 618.350000 ;
      RECT 357.500000 617.650000 383.500000 618.350000 ;
      RECT 1157.500000 616.350000 1158.500000 617.650000 ;
      RECT 1139.000000 616.350000 1149.500000 619.650000 ;
      RECT 396.500000 616.350000 399.000000 619.650000 ;
      RECT 382.500000 616.350000 383.500000 617.650000 ;
      RECT 357.500000 616.350000 358.500000 617.650000 ;
      RECT 0.000000 616.350000 349.500000 619.650000 ;
      RECT 1139.000000 615.650000 1158.500000 616.350000 ;
      RECT 382.500000 615.650000 399.000000 616.350000 ;
      RECT 0.000000 615.650000 358.500000 616.350000 ;
      RECT 1166.500000 614.350000 1186.000000 617.650000 ;
      RECT 1157.500000 614.350000 1158.500000 615.650000 ;
      RECT 382.500000 614.350000 383.500000 615.650000 ;
      RECT 366.500000 614.350000 369.500000 617.650000 ;
      RECT 357.500000 614.350000 358.500000 615.650000 ;
      RECT 1157.500000 613.650000 1186.000000 614.350000 ;
      RECT 357.500000 613.650000 383.500000 614.350000 ;
      RECT 1157.500000 612.350000 1158.500000 613.650000 ;
      RECT 1139.000000 612.350000 1149.500000 615.650000 ;
      RECT 396.500000 612.350000 399.000000 615.650000 ;
      RECT 382.500000 612.350000 383.500000 613.650000 ;
      RECT 357.500000 612.350000 358.500000 613.650000 ;
      RECT 0.000000 612.350000 349.500000 615.650000 ;
      RECT 1139.000000 611.650000 1158.500000 612.350000 ;
      RECT 382.500000 611.650000 399.000000 612.350000 ;
      RECT 0.000000 611.650000 358.500000 612.350000 ;
      RECT 1166.500000 610.350000 1186.000000 613.650000 ;
      RECT 1157.500000 610.350000 1158.500000 611.650000 ;
      RECT 382.500000 610.350000 383.500000 611.650000 ;
      RECT 366.500000 610.350000 369.500000 613.650000 ;
      RECT 357.500000 610.350000 358.500000 611.650000 ;
      RECT 1157.500000 609.650000 1186.000000 610.350000 ;
      RECT 357.500000 609.650000 383.500000 610.350000 ;
      RECT 1157.500000 608.350000 1158.500000 609.650000 ;
      RECT 1139.000000 608.350000 1149.500000 611.650000 ;
      RECT 396.500000 608.350000 399.000000 611.650000 ;
      RECT 382.500000 608.350000 383.500000 609.650000 ;
      RECT 357.500000 608.350000 358.500000 609.650000 ;
      RECT 0.000000 608.350000 349.500000 611.650000 ;
      RECT 1139.000000 607.650000 1158.500000 608.350000 ;
      RECT 382.500000 607.650000 399.000000 608.350000 ;
      RECT 0.000000 607.650000 358.500000 608.350000 ;
      RECT 1166.500000 606.350000 1186.000000 609.650000 ;
      RECT 1157.500000 606.350000 1158.500000 607.650000 ;
      RECT 382.500000 606.350000 383.500000 607.650000 ;
      RECT 366.500000 606.350000 369.500000 609.650000 ;
      RECT 357.500000 606.350000 358.500000 607.650000 ;
      RECT 1157.500000 605.650000 1186.000000 606.350000 ;
      RECT 357.500000 605.650000 383.500000 606.350000 ;
      RECT 1157.500000 604.350000 1158.500000 605.650000 ;
      RECT 1139.000000 604.350000 1149.500000 607.650000 ;
      RECT 396.500000 604.350000 399.000000 607.650000 ;
      RECT 382.500000 604.350000 383.500000 605.650000 ;
      RECT 357.500000 604.350000 358.500000 605.650000 ;
      RECT 0.000000 604.350000 349.500000 607.650000 ;
      RECT 1139.000000 603.650000 1158.500000 604.350000 ;
      RECT 382.500000 603.650000 399.000000 604.350000 ;
      RECT 0.000000 603.650000 358.500000 604.350000 ;
      RECT 1166.500000 602.350000 1186.000000 605.650000 ;
      RECT 1157.500000 602.350000 1158.500000 603.650000 ;
      RECT 382.500000 602.350000 383.500000 603.650000 ;
      RECT 366.500000 602.350000 369.500000 605.650000 ;
      RECT 357.500000 602.350000 358.500000 603.650000 ;
      RECT 1157.500000 601.650000 1186.000000 602.350000 ;
      RECT 357.500000 601.650000 383.500000 602.350000 ;
      RECT 1157.500000 600.350000 1158.500000 601.650000 ;
      RECT 1139.000000 600.350000 1149.500000 603.650000 ;
      RECT 396.500000 600.350000 399.000000 603.650000 ;
      RECT 382.500000 600.350000 383.500000 601.650000 ;
      RECT 357.500000 600.350000 358.500000 601.650000 ;
      RECT 0.000000 600.350000 349.500000 603.650000 ;
      RECT 1139.000000 599.650000 1158.500000 600.350000 ;
      RECT 382.500000 599.650000 399.000000 600.350000 ;
      RECT 0.000000 599.650000 358.500000 600.350000 ;
      RECT 1166.500000 598.350000 1186.000000 601.650000 ;
      RECT 1157.500000 598.350000 1158.500000 599.650000 ;
      RECT 382.500000 598.350000 383.500000 599.650000 ;
      RECT 366.500000 598.350000 369.500000 601.650000 ;
      RECT 357.500000 598.350000 358.500000 599.650000 ;
      RECT 1157.500000 597.650000 1186.000000 598.350000 ;
      RECT 357.500000 597.650000 383.500000 598.350000 ;
      RECT 1157.500000 596.350000 1158.500000 597.650000 ;
      RECT 1139.000000 596.350000 1149.500000 599.650000 ;
      RECT 396.500000 596.350000 399.000000 599.650000 ;
      RECT 382.500000 596.350000 383.500000 597.650000 ;
      RECT 357.500000 596.350000 358.500000 597.650000 ;
      RECT 0.000000 596.350000 349.500000 599.650000 ;
      RECT 1139.000000 595.650000 1158.500000 596.350000 ;
      RECT 382.500000 595.650000 399.000000 596.350000 ;
      RECT 0.000000 595.650000 358.500000 596.350000 ;
      RECT 1166.500000 594.350000 1186.000000 597.650000 ;
      RECT 1157.500000 594.350000 1158.500000 595.650000 ;
      RECT 382.500000 594.350000 383.500000 595.650000 ;
      RECT 366.500000 594.350000 369.500000 597.650000 ;
      RECT 357.500000 594.350000 358.500000 595.650000 ;
      RECT 1157.500000 593.650000 1186.000000 594.350000 ;
      RECT 357.500000 593.650000 383.500000 594.350000 ;
      RECT 1157.500000 592.350000 1158.500000 593.650000 ;
      RECT 1139.000000 592.350000 1149.500000 595.650000 ;
      RECT 396.500000 592.350000 399.000000 595.650000 ;
      RECT 382.500000 592.350000 383.500000 593.650000 ;
      RECT 357.500000 592.350000 358.500000 593.650000 ;
      RECT 0.000000 592.350000 349.500000 595.650000 ;
      RECT 1139.000000 591.650000 1158.500000 592.350000 ;
      RECT 382.500000 591.650000 399.000000 592.350000 ;
      RECT 0.000000 591.650000 358.500000 592.350000 ;
      RECT 1166.500000 590.350000 1186.000000 593.650000 ;
      RECT 1157.500000 590.350000 1158.500000 591.650000 ;
      RECT 382.500000 590.350000 383.500000 591.650000 ;
      RECT 366.500000 590.350000 369.500000 593.650000 ;
      RECT 357.500000 590.350000 358.500000 591.650000 ;
      RECT 1157.500000 589.650000 1186.000000 590.350000 ;
      RECT 357.500000 589.650000 383.500000 590.350000 ;
      RECT 1157.500000 588.350000 1158.500000 589.650000 ;
      RECT 1139.000000 588.350000 1149.500000 591.650000 ;
      RECT 396.500000 588.350000 399.000000 591.650000 ;
      RECT 382.500000 588.350000 383.500000 589.650000 ;
      RECT 357.500000 588.350000 358.500000 589.650000 ;
      RECT 0.000000 588.350000 349.500000 591.650000 ;
      RECT 1139.000000 587.650000 1158.500000 588.350000 ;
      RECT 382.500000 587.650000 399.000000 588.350000 ;
      RECT 0.000000 587.650000 358.500000 588.350000 ;
      RECT 1166.500000 586.350000 1186.000000 589.650000 ;
      RECT 1157.500000 586.350000 1158.500000 587.650000 ;
      RECT 382.500000 586.350000 383.500000 587.650000 ;
      RECT 366.500000 586.350000 369.500000 589.650000 ;
      RECT 357.500000 586.350000 358.500000 587.650000 ;
      RECT 1157.500000 585.650000 1186.000000 586.350000 ;
      RECT 357.500000 585.650000 383.500000 586.350000 ;
      RECT 1157.500000 584.350000 1158.500000 585.650000 ;
      RECT 1139.000000 584.350000 1149.500000 587.650000 ;
      RECT 396.500000 584.350000 399.000000 587.650000 ;
      RECT 382.500000 584.350000 383.500000 585.650000 ;
      RECT 357.500000 584.350000 358.500000 585.650000 ;
      RECT 0.000000 584.350000 349.500000 587.650000 ;
      RECT 1139.000000 583.650000 1158.500000 584.350000 ;
      RECT 382.500000 583.650000 399.000000 584.350000 ;
      RECT 0.000000 583.650000 358.500000 584.350000 ;
      RECT 1166.500000 582.350000 1186.000000 585.650000 ;
      RECT 1157.500000 582.350000 1158.500000 583.650000 ;
      RECT 382.500000 582.350000 383.500000 583.650000 ;
      RECT 366.500000 582.350000 369.500000 585.650000 ;
      RECT 357.500000 582.350000 358.500000 583.650000 ;
      RECT 1157.500000 581.650000 1186.000000 582.350000 ;
      RECT 357.500000 581.650000 383.500000 582.350000 ;
      RECT 1157.500000 580.350000 1158.500000 581.650000 ;
      RECT 1139.000000 580.350000 1149.500000 583.650000 ;
      RECT 396.500000 580.350000 399.000000 583.650000 ;
      RECT 382.500000 580.350000 383.500000 581.650000 ;
      RECT 357.500000 580.350000 358.500000 581.650000 ;
      RECT 0.000000 580.350000 349.500000 583.650000 ;
      RECT 1139.000000 579.650000 1158.500000 580.350000 ;
      RECT 382.500000 579.650000 399.000000 580.350000 ;
      RECT 0.000000 579.650000 358.500000 580.350000 ;
      RECT 1166.500000 578.350000 1186.000000 581.650000 ;
      RECT 1157.500000 578.350000 1158.500000 579.650000 ;
      RECT 382.500000 578.350000 383.500000 579.650000 ;
      RECT 366.500000 578.350000 369.500000 581.650000 ;
      RECT 357.500000 578.350000 358.500000 579.650000 ;
      RECT 1157.500000 577.650000 1186.000000 578.350000 ;
      RECT 357.500000 577.650000 383.500000 578.350000 ;
      RECT 1157.500000 576.350000 1158.500000 577.650000 ;
      RECT 1139.000000 576.350000 1149.500000 579.650000 ;
      RECT 396.500000 576.350000 399.000000 579.650000 ;
      RECT 382.500000 576.350000 383.500000 577.650000 ;
      RECT 357.500000 576.350000 358.500000 577.650000 ;
      RECT 0.000000 576.350000 349.500000 579.650000 ;
      RECT 1139.000000 575.650000 1158.500000 576.350000 ;
      RECT 382.500000 575.650000 399.000000 576.350000 ;
      RECT 0.000000 575.650000 358.500000 576.350000 ;
      RECT 1166.500000 574.350000 1186.000000 577.650000 ;
      RECT 1157.500000 574.350000 1158.500000 575.650000 ;
      RECT 382.500000 574.350000 383.500000 575.650000 ;
      RECT 366.500000 574.350000 369.500000 577.650000 ;
      RECT 357.500000 574.350000 358.500000 575.650000 ;
      RECT 1157.500000 573.650000 1186.000000 574.350000 ;
      RECT 357.500000 573.650000 383.500000 574.350000 ;
      RECT 1157.500000 572.350000 1158.500000 573.650000 ;
      RECT 1139.000000 572.350000 1149.500000 575.650000 ;
      RECT 396.500000 572.350000 399.000000 575.650000 ;
      RECT 382.500000 572.350000 383.500000 573.650000 ;
      RECT 357.500000 572.350000 358.500000 573.650000 ;
      RECT 0.000000 572.350000 349.500000 575.650000 ;
      RECT 1139.000000 571.650000 1158.500000 572.350000 ;
      RECT 382.500000 571.650000 399.000000 572.350000 ;
      RECT 0.000000 571.650000 358.500000 572.350000 ;
      RECT 1166.500000 570.350000 1186.000000 573.650000 ;
      RECT 1157.500000 570.350000 1158.500000 571.650000 ;
      RECT 382.500000 570.350000 383.500000 571.650000 ;
      RECT 366.500000 570.350000 369.500000 573.650000 ;
      RECT 357.500000 570.350000 358.500000 571.650000 ;
      RECT 1157.500000 569.650000 1186.000000 570.350000 ;
      RECT 357.500000 569.650000 383.500000 570.350000 ;
      RECT 1157.500000 568.350000 1158.500000 569.650000 ;
      RECT 1139.000000 568.350000 1149.500000 571.650000 ;
      RECT 396.500000 568.350000 399.000000 571.650000 ;
      RECT 382.500000 568.350000 383.500000 569.650000 ;
      RECT 357.500000 568.350000 358.500000 569.650000 ;
      RECT 0.000000 568.350000 349.500000 571.650000 ;
      RECT 1139.000000 567.650000 1158.500000 568.350000 ;
      RECT 382.500000 567.650000 399.000000 568.350000 ;
      RECT 0.000000 567.650000 358.500000 568.350000 ;
      RECT 1166.500000 566.350000 1186.000000 569.650000 ;
      RECT 1157.500000 566.350000 1158.500000 567.650000 ;
      RECT 382.500000 566.350000 383.500000 567.650000 ;
      RECT 366.500000 566.350000 369.500000 569.650000 ;
      RECT 357.500000 566.350000 358.500000 567.650000 ;
      RECT 1157.500000 565.650000 1186.000000 566.350000 ;
      RECT 357.500000 565.650000 383.500000 566.350000 ;
      RECT 1157.500000 564.350000 1158.500000 565.650000 ;
      RECT 1139.000000 564.350000 1149.500000 567.650000 ;
      RECT 396.500000 564.350000 399.000000 567.650000 ;
      RECT 382.500000 564.350000 383.500000 565.650000 ;
      RECT 357.500000 564.350000 358.500000 565.650000 ;
      RECT 0.000000 564.350000 349.500000 567.650000 ;
      RECT 1139.000000 563.650000 1158.500000 564.350000 ;
      RECT 382.500000 563.650000 399.000000 564.350000 ;
      RECT 0.000000 563.650000 358.500000 564.350000 ;
      RECT 1166.500000 562.350000 1186.000000 565.650000 ;
      RECT 1157.500000 562.350000 1158.500000 563.650000 ;
      RECT 382.500000 562.350000 383.500000 563.650000 ;
      RECT 366.500000 562.350000 369.500000 565.650000 ;
      RECT 357.500000 562.350000 358.500000 563.650000 ;
      RECT 1157.500000 561.650000 1186.000000 562.350000 ;
      RECT 357.500000 561.650000 383.500000 562.350000 ;
      RECT 1157.500000 560.350000 1158.500000 561.650000 ;
      RECT 1139.000000 560.350000 1149.500000 563.650000 ;
      RECT 396.500000 560.350000 399.000000 563.650000 ;
      RECT 382.500000 560.350000 383.500000 561.650000 ;
      RECT 357.500000 560.350000 358.500000 561.650000 ;
      RECT 0.000000 560.350000 349.500000 563.650000 ;
      RECT 1139.000000 559.650000 1158.500000 560.350000 ;
      RECT 382.500000 559.650000 399.000000 560.350000 ;
      RECT 0.000000 559.650000 358.500000 560.350000 ;
      RECT 1166.500000 558.350000 1186.000000 561.650000 ;
      RECT 1157.500000 558.350000 1158.500000 559.650000 ;
      RECT 382.500000 558.350000 383.500000 559.650000 ;
      RECT 366.500000 558.350000 369.500000 561.650000 ;
      RECT 357.500000 558.350000 358.500000 559.650000 ;
      RECT 1157.500000 557.650000 1186.000000 558.350000 ;
      RECT 357.500000 557.650000 383.500000 558.350000 ;
      RECT 1157.500000 556.350000 1158.500000 557.650000 ;
      RECT 1139.000000 556.350000 1149.500000 559.650000 ;
      RECT 396.500000 556.350000 399.000000 559.650000 ;
      RECT 382.500000 556.350000 383.500000 557.650000 ;
      RECT 357.500000 556.350000 358.500000 557.650000 ;
      RECT 0.000000 556.350000 349.500000 559.650000 ;
      RECT 1139.000000 555.650000 1158.500000 556.350000 ;
      RECT 382.500000 555.650000 399.000000 556.350000 ;
      RECT 0.000000 555.650000 358.500000 556.350000 ;
      RECT 1166.500000 554.350000 1186.000000 557.650000 ;
      RECT 1157.500000 554.350000 1158.500000 555.650000 ;
      RECT 382.500000 554.350000 383.500000 555.650000 ;
      RECT 366.500000 554.350000 369.500000 557.650000 ;
      RECT 357.500000 554.350000 358.500000 555.650000 ;
      RECT 1157.500000 553.650000 1186.000000 554.350000 ;
      RECT 357.500000 553.650000 383.500000 554.350000 ;
      RECT 1157.500000 552.350000 1158.500000 553.650000 ;
      RECT 1139.000000 552.350000 1149.500000 555.650000 ;
      RECT 396.500000 552.350000 399.000000 555.650000 ;
      RECT 382.500000 552.350000 383.500000 553.650000 ;
      RECT 357.500000 552.350000 358.500000 553.650000 ;
      RECT 0.000000 552.350000 349.500000 555.650000 ;
      RECT 1139.000000 551.650000 1158.500000 552.350000 ;
      RECT 382.500000 551.650000 399.000000 552.350000 ;
      RECT 0.000000 551.650000 358.500000 552.350000 ;
      RECT 1166.500000 550.350000 1186.000000 553.650000 ;
      RECT 1157.500000 550.350000 1158.500000 551.650000 ;
      RECT 382.500000 550.350000 383.500000 551.650000 ;
      RECT 366.500000 550.350000 369.500000 553.650000 ;
      RECT 357.500000 550.350000 358.500000 551.650000 ;
      RECT 1157.500000 549.650000 1186.000000 550.350000 ;
      RECT 357.500000 549.650000 383.500000 550.350000 ;
      RECT 1157.500000 548.350000 1158.500000 549.650000 ;
      RECT 1139.000000 548.350000 1149.500000 551.650000 ;
      RECT 396.500000 548.350000 399.000000 551.650000 ;
      RECT 382.500000 548.350000 383.500000 549.650000 ;
      RECT 357.500000 548.350000 358.500000 549.650000 ;
      RECT 0.000000 548.350000 349.500000 551.650000 ;
      RECT 1139.000000 547.650000 1158.500000 548.350000 ;
      RECT 382.500000 547.650000 399.000000 548.350000 ;
      RECT 0.000000 547.650000 358.500000 548.350000 ;
      RECT 1166.500000 546.350000 1186.000000 549.650000 ;
      RECT 1157.500000 546.350000 1158.500000 547.650000 ;
      RECT 382.500000 546.350000 383.500000 547.650000 ;
      RECT 366.500000 546.350000 369.500000 549.650000 ;
      RECT 357.500000 546.350000 358.500000 547.650000 ;
      RECT 1157.500000 545.650000 1186.000000 546.350000 ;
      RECT 357.500000 545.650000 383.500000 546.350000 ;
      RECT 1157.500000 544.350000 1158.500000 545.650000 ;
      RECT 1139.000000 544.350000 1149.500000 547.650000 ;
      RECT 396.500000 544.350000 399.000000 547.650000 ;
      RECT 382.500000 544.350000 383.500000 545.650000 ;
      RECT 357.500000 544.350000 358.500000 545.650000 ;
      RECT 0.000000 544.350000 349.500000 547.650000 ;
      RECT 1139.000000 543.650000 1158.500000 544.350000 ;
      RECT 382.500000 543.650000 399.000000 544.350000 ;
      RECT 0.000000 543.650000 358.500000 544.350000 ;
      RECT 1166.500000 542.350000 1186.000000 545.650000 ;
      RECT 1157.500000 542.350000 1158.500000 543.650000 ;
      RECT 382.500000 542.350000 383.500000 543.650000 ;
      RECT 366.500000 542.350000 369.500000 545.650000 ;
      RECT 357.500000 542.350000 358.500000 543.650000 ;
      RECT 1157.500000 541.650000 1186.000000 542.350000 ;
      RECT 357.500000 541.650000 383.500000 542.350000 ;
      RECT 1157.500000 540.350000 1158.500000 541.650000 ;
      RECT 1139.000000 540.350000 1149.500000 543.650000 ;
      RECT 396.500000 540.350000 399.000000 543.650000 ;
      RECT 382.500000 540.350000 383.500000 541.650000 ;
      RECT 357.500000 540.350000 358.500000 541.650000 ;
      RECT 0.000000 540.350000 349.500000 543.650000 ;
      RECT 1139.000000 539.650000 1158.500000 540.350000 ;
      RECT 382.500000 539.650000 399.000000 540.350000 ;
      RECT 0.000000 539.650000 358.500000 540.350000 ;
      RECT 1166.500000 538.350000 1186.000000 541.650000 ;
      RECT 1157.500000 538.350000 1158.500000 539.650000 ;
      RECT 382.500000 538.350000 383.500000 539.650000 ;
      RECT 366.500000 538.350000 369.500000 541.650000 ;
      RECT 357.500000 538.350000 358.500000 539.650000 ;
      RECT 1157.500000 537.650000 1186.000000 538.350000 ;
      RECT 357.500000 537.650000 383.500000 538.350000 ;
      RECT 1157.500000 536.350000 1158.500000 537.650000 ;
      RECT 1139.000000 536.350000 1149.500000 539.650000 ;
      RECT 396.500000 536.350000 399.000000 539.650000 ;
      RECT 382.500000 536.350000 383.500000 537.650000 ;
      RECT 357.500000 536.350000 358.500000 537.650000 ;
      RECT 0.000000 536.350000 349.500000 539.650000 ;
      RECT 1139.000000 535.650000 1158.500000 536.350000 ;
      RECT 382.500000 535.650000 399.000000 536.350000 ;
      RECT 0.000000 535.650000 358.500000 536.350000 ;
      RECT 1166.500000 534.350000 1186.000000 537.650000 ;
      RECT 1157.500000 534.350000 1158.500000 535.650000 ;
      RECT 382.500000 534.350000 383.500000 535.650000 ;
      RECT 366.500000 534.350000 369.500000 537.650000 ;
      RECT 357.500000 534.350000 358.500000 535.650000 ;
      RECT 1157.500000 533.650000 1186.000000 534.350000 ;
      RECT 357.500000 533.650000 383.500000 534.350000 ;
      RECT 1157.500000 532.350000 1158.500000 533.650000 ;
      RECT 1139.000000 532.350000 1149.500000 535.650000 ;
      RECT 396.500000 532.350000 399.000000 535.650000 ;
      RECT 382.500000 532.350000 383.500000 533.650000 ;
      RECT 357.500000 532.350000 358.500000 533.650000 ;
      RECT 0.000000 532.350000 349.500000 535.650000 ;
      RECT 1139.000000 531.650000 1158.500000 532.350000 ;
      RECT 382.500000 531.650000 399.000000 532.350000 ;
      RECT 0.000000 531.650000 358.500000 532.350000 ;
      RECT 1166.500000 530.350000 1186.000000 533.650000 ;
      RECT 1157.500000 530.350000 1158.500000 531.650000 ;
      RECT 382.500000 530.350000 383.500000 531.650000 ;
      RECT 366.500000 530.350000 369.500000 533.650000 ;
      RECT 357.500000 530.350000 358.500000 531.650000 ;
      RECT 1157.500000 529.650000 1186.000000 530.350000 ;
      RECT 357.500000 529.650000 383.500000 530.350000 ;
      RECT 1157.500000 528.350000 1158.500000 529.650000 ;
      RECT 1139.000000 528.350000 1149.500000 531.650000 ;
      RECT 396.500000 528.350000 399.000000 531.650000 ;
      RECT 382.500000 528.350000 383.500000 529.650000 ;
      RECT 357.500000 528.350000 358.500000 529.650000 ;
      RECT 0.000000 528.350000 349.500000 531.650000 ;
      RECT 1139.000000 527.650000 1158.500000 528.350000 ;
      RECT 382.500000 527.650000 399.000000 528.350000 ;
      RECT 0.000000 527.650000 358.500000 528.350000 ;
      RECT 1166.500000 526.350000 1186.000000 529.650000 ;
      RECT 1157.500000 526.350000 1158.500000 527.650000 ;
      RECT 382.500000 526.350000 383.500000 527.650000 ;
      RECT 366.500000 526.350000 369.500000 529.650000 ;
      RECT 357.500000 526.350000 358.500000 527.650000 ;
      RECT 1157.500000 525.650000 1186.000000 526.350000 ;
      RECT 357.500000 525.650000 383.500000 526.350000 ;
      RECT 1157.500000 524.350000 1158.500000 525.650000 ;
      RECT 1139.000000 524.350000 1149.500000 527.650000 ;
      RECT 396.500000 524.350000 399.000000 527.650000 ;
      RECT 382.500000 524.350000 383.500000 525.650000 ;
      RECT 357.500000 524.350000 358.500000 525.650000 ;
      RECT 0.000000 524.350000 349.500000 527.650000 ;
      RECT 1139.000000 523.650000 1158.500000 524.350000 ;
      RECT 382.500000 523.650000 399.000000 524.350000 ;
      RECT 0.000000 523.650000 358.500000 524.350000 ;
      RECT 1166.500000 522.350000 1186.000000 525.650000 ;
      RECT 1157.500000 522.350000 1158.500000 523.650000 ;
      RECT 382.500000 522.350000 383.500000 523.650000 ;
      RECT 366.500000 522.350000 369.500000 525.650000 ;
      RECT 357.500000 522.350000 358.500000 523.650000 ;
      RECT 1157.500000 521.650000 1186.000000 522.350000 ;
      RECT 357.500000 521.650000 383.500000 522.350000 ;
      RECT 1157.500000 520.350000 1158.500000 521.650000 ;
      RECT 1139.000000 520.350000 1149.500000 523.650000 ;
      RECT 396.500000 520.350000 399.000000 523.650000 ;
      RECT 382.500000 520.350000 383.500000 521.650000 ;
      RECT 357.500000 520.350000 358.500000 521.650000 ;
      RECT 0.000000 520.350000 349.500000 523.650000 ;
      RECT 1139.000000 519.650000 1158.500000 520.350000 ;
      RECT 382.500000 519.650000 399.000000 520.350000 ;
      RECT 0.000000 519.650000 358.500000 520.350000 ;
      RECT 1166.500000 518.350000 1186.000000 521.650000 ;
      RECT 1157.500000 518.350000 1158.500000 519.650000 ;
      RECT 382.500000 518.350000 383.500000 519.650000 ;
      RECT 366.500000 518.350000 369.500000 521.650000 ;
      RECT 357.500000 518.350000 358.500000 519.650000 ;
      RECT 1157.500000 517.650000 1186.000000 518.350000 ;
      RECT 357.500000 517.650000 383.500000 518.350000 ;
      RECT 307.500000 517.650000 349.500000 519.650000 ;
      RECT 0.000000 517.650000 299.500000 519.650000 ;
      RECT 1157.500000 516.350000 1158.500000 517.650000 ;
      RECT 1139.000000 516.350000 1149.500000 519.650000 ;
      RECT 396.500000 516.350000 399.000000 519.650000 ;
      RECT 382.500000 516.350000 383.500000 517.650000 ;
      RECT 357.500000 516.350000 358.500000 517.650000 ;
      RECT 316.500000 516.350000 349.500000 517.650000 ;
      RECT 307.500000 516.350000 308.500000 517.650000 ;
      RECT 266.500000 516.350000 299.500000 517.650000 ;
      RECT 1139.000000 515.650000 1158.500000 516.350000 ;
      RECT 382.500000 515.650000 399.000000 516.350000 ;
      RECT 316.500000 515.650000 358.500000 516.350000 ;
      RECT 266.500000 515.650000 308.500000 516.350000 ;
      RECT 216.500000 515.650000 258.500000 517.650000 ;
      RECT 166.500000 515.650000 208.500000 517.650000 ;
      RECT 116.500000 515.650000 158.500000 517.650000 ;
      RECT 66.500000 515.650000 108.500000 517.650000 ;
      RECT 29.500000 515.650000 58.500000 517.650000 ;
      RECT 0.000000 515.650000 16.500000 517.650000 ;
      RECT 1166.500000 514.350000 1186.000000 517.650000 ;
      RECT 1157.500000 514.350000 1158.500000 515.650000 ;
      RECT 382.500000 514.350000 383.500000 515.650000 ;
      RECT 366.500000 514.350000 369.500000 517.650000 ;
      RECT 357.500000 514.350000 358.500000 515.650000 ;
      RECT 316.500000 514.350000 349.500000 515.650000 ;
      RECT 307.500000 514.350000 308.500000 515.650000 ;
      RECT 266.500000 514.350000 299.500000 515.650000 ;
      RECT 257.500000 514.350000 258.500000 515.650000 ;
      RECT 216.500000 514.350000 249.500000 515.650000 ;
      RECT 207.500000 514.350000 208.500000 515.650000 ;
      RECT 166.500000 514.350000 199.500000 515.650000 ;
      RECT 157.500000 514.350000 158.500000 515.650000 ;
      RECT 116.500000 514.350000 149.500000 515.650000 ;
      RECT 107.500000 514.350000 108.500000 515.650000 ;
      RECT 66.500000 514.350000 99.500000 515.650000 ;
      RECT 57.500000 514.350000 58.500000 515.650000 ;
      RECT 29.500000 514.350000 49.500000 515.650000 ;
      RECT 15.500000 514.350000 16.500000 515.650000 ;
      RECT 1157.500000 513.650000 1186.000000 514.350000 ;
      RECT 357.500000 513.650000 383.500000 514.350000 ;
      RECT 307.500000 513.650000 349.500000 514.350000 ;
      RECT 257.500000 513.650000 299.500000 514.350000 ;
      RECT 207.500000 513.650000 249.500000 514.350000 ;
      RECT 157.500000 513.650000 199.500000 514.350000 ;
      RECT 107.500000 513.650000 149.500000 514.350000 ;
      RECT 57.500000 513.650000 99.500000 514.350000 ;
      RECT 15.500000 513.650000 49.500000 514.350000 ;
      RECT 1157.500000 512.350000 1158.500000 513.650000 ;
      RECT 1139.000000 512.350000 1149.500000 515.650000 ;
      RECT 396.500000 512.350000 399.000000 515.650000 ;
      RECT 382.500000 512.350000 383.500000 513.650000 ;
      RECT 357.500000 512.350000 358.500000 513.650000 ;
      RECT 316.500000 512.350000 349.500000 513.650000 ;
      RECT 307.500000 512.350000 308.500000 513.650000 ;
      RECT 266.500000 512.350000 299.500000 513.650000 ;
      RECT 257.500000 512.350000 258.500000 513.650000 ;
      RECT 216.500000 512.350000 249.500000 513.650000 ;
      RECT 207.500000 512.350000 208.500000 513.650000 ;
      RECT 166.500000 512.350000 199.500000 513.650000 ;
      RECT 157.500000 512.350000 158.500000 513.650000 ;
      RECT 116.500000 512.350000 149.500000 513.650000 ;
      RECT 107.500000 512.350000 108.500000 513.650000 ;
      RECT 66.500000 512.350000 99.500000 513.650000 ;
      RECT 57.500000 512.350000 58.500000 513.650000 ;
      RECT 29.500000 512.350000 49.500000 513.650000 ;
      RECT 15.500000 512.350000 16.500000 513.650000 ;
      RECT 0.000000 512.350000 2.500000 515.650000 ;
      RECT 1139.000000 511.650000 1158.500000 512.350000 ;
      RECT 382.500000 511.650000 399.000000 512.350000 ;
      RECT 316.500000 511.650000 358.500000 512.350000 ;
      RECT 266.500000 511.650000 308.500000 512.350000 ;
      RECT 216.500000 511.650000 258.500000 512.350000 ;
      RECT 166.500000 511.650000 208.500000 512.350000 ;
      RECT 116.500000 511.650000 158.500000 512.350000 ;
      RECT 66.500000 511.650000 108.500000 512.350000 ;
      RECT 29.500000 511.650000 58.500000 512.350000 ;
      RECT 0.000000 511.650000 16.500000 512.350000 ;
      RECT 1166.500000 510.350000 1186.000000 513.650000 ;
      RECT 1157.500000 510.350000 1158.500000 511.650000 ;
      RECT 382.500000 510.350000 383.500000 511.650000 ;
      RECT 366.500000 510.350000 369.500000 513.650000 ;
      RECT 357.500000 510.350000 358.500000 511.650000 ;
      RECT 316.500000 510.350000 349.500000 511.650000 ;
      RECT 307.500000 510.350000 308.500000 511.650000 ;
      RECT 266.500000 510.350000 299.500000 511.650000 ;
      RECT 257.500000 510.350000 258.500000 511.650000 ;
      RECT 216.500000 510.350000 249.500000 511.650000 ;
      RECT 207.500000 510.350000 208.500000 511.650000 ;
      RECT 166.500000 510.350000 199.500000 511.650000 ;
      RECT 157.500000 510.350000 158.500000 511.650000 ;
      RECT 116.500000 510.350000 149.500000 511.650000 ;
      RECT 107.500000 510.350000 108.500000 511.650000 ;
      RECT 66.500000 510.350000 99.500000 511.650000 ;
      RECT 57.500000 510.350000 58.500000 511.650000 ;
      RECT 29.500000 510.350000 49.500000 511.650000 ;
      RECT 15.500000 510.350000 16.500000 511.650000 ;
      RECT 1157.500000 509.650000 1186.000000 510.350000 ;
      RECT 357.500000 509.650000 383.500000 510.350000 ;
      RECT 307.500000 509.650000 349.500000 510.350000 ;
      RECT 257.500000 509.650000 299.500000 510.350000 ;
      RECT 207.500000 509.650000 249.500000 510.350000 ;
      RECT 157.500000 509.650000 199.500000 510.350000 ;
      RECT 107.500000 509.650000 149.500000 510.350000 ;
      RECT 57.500000 509.650000 99.500000 510.350000 ;
      RECT 15.500000 509.650000 49.500000 510.350000 ;
      RECT 1157.500000 508.350000 1158.500000 509.650000 ;
      RECT 1139.000000 508.350000 1149.500000 511.650000 ;
      RECT 396.500000 508.350000 399.000000 511.650000 ;
      RECT 382.500000 508.350000 383.500000 509.650000 ;
      RECT 357.500000 508.350000 358.500000 509.650000 ;
      RECT 316.500000 508.350000 349.500000 509.650000 ;
      RECT 307.500000 508.350000 308.500000 509.650000 ;
      RECT 266.500000 508.350000 299.500000 509.650000 ;
      RECT 257.500000 508.350000 258.500000 509.650000 ;
      RECT 216.500000 508.350000 249.500000 509.650000 ;
      RECT 207.500000 508.350000 208.500000 509.650000 ;
      RECT 166.500000 508.350000 199.500000 509.650000 ;
      RECT 157.500000 508.350000 158.500000 509.650000 ;
      RECT 116.500000 508.350000 149.500000 509.650000 ;
      RECT 107.500000 508.350000 108.500000 509.650000 ;
      RECT 66.500000 508.350000 99.500000 509.650000 ;
      RECT 57.500000 508.350000 58.500000 509.650000 ;
      RECT 29.500000 508.350000 49.500000 509.650000 ;
      RECT 15.500000 508.350000 16.500000 509.650000 ;
      RECT 0.000000 508.350000 2.500000 511.650000 ;
      RECT 1139.000000 507.650000 1158.500000 508.350000 ;
      RECT 382.500000 507.650000 399.000000 508.350000 ;
      RECT 316.500000 507.650000 358.500000 508.350000 ;
      RECT 266.500000 507.650000 308.500000 508.350000 ;
      RECT 216.500000 507.650000 258.500000 508.350000 ;
      RECT 166.500000 507.650000 208.500000 508.350000 ;
      RECT 116.500000 507.650000 158.500000 508.350000 ;
      RECT 66.500000 507.650000 108.500000 508.350000 ;
      RECT 29.500000 507.650000 58.500000 508.350000 ;
      RECT 0.000000 507.650000 16.500000 508.350000 ;
      RECT 1166.500000 506.350000 1186.000000 509.650000 ;
      RECT 1157.500000 506.350000 1158.500000 507.650000 ;
      RECT 382.500000 506.350000 383.500000 507.650000 ;
      RECT 366.500000 506.350000 369.500000 509.650000 ;
      RECT 357.500000 506.350000 358.500000 507.650000 ;
      RECT 316.500000 506.350000 349.500000 507.650000 ;
      RECT 307.500000 506.350000 308.500000 507.650000 ;
      RECT 266.500000 506.350000 299.500000 507.650000 ;
      RECT 257.500000 506.350000 258.500000 507.650000 ;
      RECT 216.500000 506.350000 249.500000 507.650000 ;
      RECT 207.500000 506.350000 208.500000 507.650000 ;
      RECT 166.500000 506.350000 199.500000 507.650000 ;
      RECT 157.500000 506.350000 158.500000 507.650000 ;
      RECT 116.500000 506.350000 149.500000 507.650000 ;
      RECT 107.500000 506.350000 108.500000 507.650000 ;
      RECT 66.500000 506.350000 99.500000 507.650000 ;
      RECT 57.500000 506.350000 58.500000 507.650000 ;
      RECT 29.500000 506.350000 49.500000 507.650000 ;
      RECT 15.500000 506.350000 16.500000 507.650000 ;
      RECT 396.500000 506.000000 399.000000 507.650000 ;
      RECT 1157.500000 505.650000 1186.000000 506.350000 ;
      RECT 396.500000 505.650000 749.000000 506.000000 ;
      RECT 357.500000 505.650000 383.500000 506.350000 ;
      RECT 307.500000 505.650000 349.500000 506.350000 ;
      RECT 257.500000 505.650000 299.500000 506.350000 ;
      RECT 207.500000 505.650000 249.500000 506.350000 ;
      RECT 157.500000 505.650000 199.500000 506.350000 ;
      RECT 107.500000 505.650000 149.500000 506.350000 ;
      RECT 57.500000 505.650000 99.500000 506.350000 ;
      RECT 15.500000 505.650000 49.500000 506.350000 ;
      RECT 1157.500000 504.350000 1158.500000 505.650000 ;
      RECT 1139.000000 504.350000 1149.500000 507.650000 ;
      RECT 396.500000 504.350000 408.500000 505.650000 ;
      RECT 382.500000 504.350000 383.500000 505.650000 ;
      RECT 357.500000 504.350000 358.500000 505.650000 ;
      RECT 316.500000 504.350000 349.500000 505.650000 ;
      RECT 307.500000 504.350000 308.500000 505.650000 ;
      RECT 266.500000 504.350000 299.500000 505.650000 ;
      RECT 257.500000 504.350000 258.500000 505.650000 ;
      RECT 216.500000 504.350000 249.500000 505.650000 ;
      RECT 207.500000 504.350000 208.500000 505.650000 ;
      RECT 166.500000 504.350000 199.500000 505.650000 ;
      RECT 157.500000 504.350000 158.500000 505.650000 ;
      RECT 116.500000 504.350000 149.500000 505.650000 ;
      RECT 107.500000 504.350000 108.500000 505.650000 ;
      RECT 66.500000 504.350000 99.500000 505.650000 ;
      RECT 57.500000 504.350000 58.500000 505.650000 ;
      RECT 29.500000 504.350000 49.500000 505.650000 ;
      RECT 15.500000 504.350000 16.500000 505.650000 ;
      RECT 0.000000 504.350000 2.500000 507.650000 ;
      RECT 1139.000000 503.650000 1158.500000 504.350000 ;
      RECT 716.500000 503.650000 749.000000 505.650000 ;
      RECT 666.500000 503.650000 708.500000 505.650000 ;
      RECT 616.500000 503.650000 658.500000 505.650000 ;
      RECT 566.500000 503.650000 608.500000 505.650000 ;
      RECT 516.500000 503.650000 558.500000 505.650000 ;
      RECT 466.500000 503.650000 508.500000 505.650000 ;
      RECT 416.500000 503.650000 458.500000 505.650000 ;
      RECT 382.500000 503.650000 408.500000 504.350000 ;
      RECT 316.500000 503.650000 358.500000 504.350000 ;
      RECT 266.500000 503.650000 308.500000 504.350000 ;
      RECT 216.500000 503.650000 258.500000 504.350000 ;
      RECT 166.500000 503.650000 208.500000 504.350000 ;
      RECT 116.500000 503.650000 158.500000 504.350000 ;
      RECT 66.500000 503.650000 108.500000 504.350000 ;
      RECT 29.500000 503.650000 58.500000 504.350000 ;
      RECT 0.000000 503.650000 16.500000 504.350000 ;
      RECT 1166.500000 502.350000 1186.000000 505.650000 ;
      RECT 1157.500000 502.350000 1158.500000 503.650000 ;
      RECT 716.500000 502.350000 733.500000 503.650000 ;
      RECT 707.500000 502.350000 708.500000 503.650000 ;
      RECT 666.500000 502.350000 699.500000 503.650000 ;
      RECT 657.500000 502.350000 658.500000 503.650000 ;
      RECT 616.500000 502.350000 649.500000 503.650000 ;
      RECT 607.500000 502.350000 608.500000 503.650000 ;
      RECT 566.500000 502.350000 599.500000 503.650000 ;
      RECT 557.500000 502.350000 558.500000 503.650000 ;
      RECT 516.500000 502.350000 549.500000 503.650000 ;
      RECT 507.500000 502.350000 508.500000 503.650000 ;
      RECT 466.500000 502.350000 499.500000 503.650000 ;
      RECT 457.500000 502.350000 458.500000 503.650000 ;
      RECT 416.500000 502.350000 449.500000 503.650000 ;
      RECT 407.500000 502.350000 408.500000 503.650000 ;
      RECT 382.500000 502.350000 383.500000 503.650000 ;
      RECT 366.500000 502.350000 369.500000 505.650000 ;
      RECT 357.500000 502.350000 358.500000 503.650000 ;
      RECT 316.500000 502.350000 349.500000 503.650000 ;
      RECT 307.500000 502.350000 308.500000 503.650000 ;
      RECT 266.500000 502.350000 299.500000 503.650000 ;
      RECT 257.500000 502.350000 258.500000 503.650000 ;
      RECT 216.500000 502.350000 249.500000 503.650000 ;
      RECT 207.500000 502.350000 208.500000 503.650000 ;
      RECT 166.500000 502.350000 199.500000 503.650000 ;
      RECT 157.500000 502.350000 158.500000 503.650000 ;
      RECT 116.500000 502.350000 149.500000 503.650000 ;
      RECT 107.500000 502.350000 108.500000 503.650000 ;
      RECT 66.500000 502.350000 99.500000 503.650000 ;
      RECT 57.500000 502.350000 58.500000 503.650000 ;
      RECT 29.500000 502.350000 49.500000 503.650000 ;
      RECT 15.500000 502.350000 16.500000 503.650000 ;
      RECT 1157.500000 501.650000 1186.000000 502.350000 ;
      RECT 707.500000 501.650000 733.500000 502.350000 ;
      RECT 657.500000 501.650000 699.500000 502.350000 ;
      RECT 607.500000 501.650000 649.500000 502.350000 ;
      RECT 557.500000 501.650000 599.500000 502.350000 ;
      RECT 507.500000 501.650000 549.500000 502.350000 ;
      RECT 457.500000 501.650000 499.500000 502.350000 ;
      RECT 407.500000 501.650000 449.500000 502.350000 ;
      RECT 357.500000 501.650000 383.500000 502.350000 ;
      RECT 307.500000 501.650000 349.500000 502.350000 ;
      RECT 257.500000 501.650000 299.500000 502.350000 ;
      RECT 207.500000 501.650000 249.500000 502.350000 ;
      RECT 157.500000 501.650000 199.500000 502.350000 ;
      RECT 107.500000 501.650000 149.500000 502.350000 ;
      RECT 57.500000 501.650000 99.500000 502.350000 ;
      RECT 15.500000 501.650000 49.500000 502.350000 ;
      RECT 1157.500000 500.350000 1158.500000 501.650000 ;
      RECT 1139.000000 500.350000 1149.500000 503.650000 ;
      RECT 746.500000 500.350000 749.000000 503.650000 ;
      RECT 716.500000 500.350000 733.500000 501.650000 ;
      RECT 707.500000 500.350000 708.500000 501.650000 ;
      RECT 666.500000 500.350000 699.500000 501.650000 ;
      RECT 657.500000 500.350000 658.500000 501.650000 ;
      RECT 616.500000 500.350000 649.500000 501.650000 ;
      RECT 607.500000 500.350000 608.500000 501.650000 ;
      RECT 566.500000 500.350000 599.500000 501.650000 ;
      RECT 557.500000 500.350000 558.500000 501.650000 ;
      RECT 516.500000 500.350000 549.500000 501.650000 ;
      RECT 507.500000 500.350000 508.500000 501.650000 ;
      RECT 466.500000 500.350000 499.500000 501.650000 ;
      RECT 457.500000 500.350000 458.500000 501.650000 ;
      RECT 416.500000 500.350000 449.500000 501.650000 ;
      RECT 407.500000 500.350000 408.500000 501.650000 ;
      RECT 396.500000 500.350000 399.500000 503.650000 ;
      RECT 382.500000 500.350000 383.500000 501.650000 ;
      RECT 357.500000 500.350000 358.500000 501.650000 ;
      RECT 316.500000 500.350000 349.500000 501.650000 ;
      RECT 307.500000 500.350000 308.500000 501.650000 ;
      RECT 266.500000 500.350000 299.500000 501.650000 ;
      RECT 257.500000 500.350000 258.500000 501.650000 ;
      RECT 216.500000 500.350000 249.500000 501.650000 ;
      RECT 207.500000 500.350000 208.500000 501.650000 ;
      RECT 166.500000 500.350000 199.500000 501.650000 ;
      RECT 157.500000 500.350000 158.500000 501.650000 ;
      RECT 116.500000 500.350000 149.500000 501.650000 ;
      RECT 107.500000 500.350000 108.500000 501.650000 ;
      RECT 66.500000 500.350000 99.500000 501.650000 ;
      RECT 57.500000 500.350000 58.500000 501.650000 ;
      RECT 29.500000 500.350000 49.500000 501.650000 ;
      RECT 15.500000 500.350000 16.500000 501.650000 ;
      RECT 0.000000 500.350000 2.500000 503.650000 ;
      RECT 1139.000000 499.650000 1158.500000 500.350000 ;
      RECT 716.500000 499.650000 749.000000 500.350000 ;
      RECT 666.500000 499.650000 708.500000 500.350000 ;
      RECT 616.500000 499.650000 658.500000 500.350000 ;
      RECT 566.500000 499.650000 608.500000 500.350000 ;
      RECT 516.500000 499.650000 558.500000 500.350000 ;
      RECT 466.500000 499.650000 508.500000 500.350000 ;
      RECT 416.500000 499.650000 458.500000 500.350000 ;
      RECT 382.500000 499.650000 408.500000 500.350000 ;
      RECT 316.500000 499.650000 358.500000 500.350000 ;
      RECT 266.500000 499.650000 308.500000 500.350000 ;
      RECT 216.500000 499.650000 258.500000 500.350000 ;
      RECT 166.500000 499.650000 208.500000 500.350000 ;
      RECT 116.500000 499.650000 158.500000 500.350000 ;
      RECT 66.500000 499.650000 108.500000 500.350000 ;
      RECT 29.500000 499.650000 58.500000 500.350000 ;
      RECT 0.000000 499.650000 16.500000 500.350000 ;
      RECT 1166.500000 498.350000 1186.000000 501.650000 ;
      RECT 1157.500000 498.350000 1158.500000 499.650000 ;
      RECT 716.500000 498.350000 733.500000 499.650000 ;
      RECT 707.500000 498.350000 708.500000 499.650000 ;
      RECT 666.500000 498.350000 699.500000 499.650000 ;
      RECT 657.500000 498.350000 658.500000 499.650000 ;
      RECT 616.500000 498.350000 649.500000 499.650000 ;
      RECT 607.500000 498.350000 608.500000 499.650000 ;
      RECT 566.500000 498.350000 599.500000 499.650000 ;
      RECT 557.500000 498.350000 558.500000 499.650000 ;
      RECT 516.500000 498.350000 549.500000 499.650000 ;
      RECT 507.500000 498.350000 508.500000 499.650000 ;
      RECT 466.500000 498.350000 499.500000 499.650000 ;
      RECT 457.500000 498.350000 458.500000 499.650000 ;
      RECT 416.500000 498.350000 449.500000 499.650000 ;
      RECT 407.500000 498.350000 408.500000 499.650000 ;
      RECT 382.500000 498.350000 383.500000 499.650000 ;
      RECT 366.500000 498.350000 369.500000 501.650000 ;
      RECT 357.500000 498.350000 358.500000 499.650000 ;
      RECT 316.500000 498.350000 349.500000 499.650000 ;
      RECT 307.500000 498.350000 308.500000 499.650000 ;
      RECT 266.500000 498.350000 299.500000 499.650000 ;
      RECT 257.500000 498.350000 258.500000 499.650000 ;
      RECT 216.500000 498.350000 249.500000 499.650000 ;
      RECT 207.500000 498.350000 208.500000 499.650000 ;
      RECT 166.500000 498.350000 199.500000 499.650000 ;
      RECT 157.500000 498.350000 158.500000 499.650000 ;
      RECT 116.500000 498.350000 149.500000 499.650000 ;
      RECT 107.500000 498.350000 108.500000 499.650000 ;
      RECT 66.500000 498.350000 99.500000 499.650000 ;
      RECT 57.500000 498.350000 58.500000 499.650000 ;
      RECT 29.500000 498.350000 49.500000 499.650000 ;
      RECT 15.500000 498.350000 16.500000 499.650000 ;
      RECT 1157.500000 497.650000 1186.000000 498.350000 ;
      RECT 707.500000 497.650000 733.500000 498.350000 ;
      RECT 657.500000 497.650000 699.500000 498.350000 ;
      RECT 607.500000 497.650000 649.500000 498.350000 ;
      RECT 557.500000 497.650000 599.500000 498.350000 ;
      RECT 507.500000 497.650000 549.500000 498.350000 ;
      RECT 457.500000 497.650000 499.500000 498.350000 ;
      RECT 407.500000 497.650000 449.500000 498.350000 ;
      RECT 357.500000 497.650000 383.500000 498.350000 ;
      RECT 307.500000 497.650000 349.500000 498.350000 ;
      RECT 257.500000 497.650000 299.500000 498.350000 ;
      RECT 207.500000 497.650000 249.500000 498.350000 ;
      RECT 157.500000 497.650000 199.500000 498.350000 ;
      RECT 107.500000 497.650000 149.500000 498.350000 ;
      RECT 57.500000 497.650000 99.500000 498.350000 ;
      RECT 15.500000 497.650000 49.500000 498.350000 ;
      RECT 1157.500000 496.350000 1158.500000 497.650000 ;
      RECT 1139.000000 496.350000 1149.500000 499.650000 ;
      RECT 746.500000 496.350000 749.000000 499.650000 ;
      RECT 716.500000 496.350000 733.500000 497.650000 ;
      RECT 707.500000 496.350000 708.500000 497.650000 ;
      RECT 666.500000 496.350000 699.500000 497.650000 ;
      RECT 657.500000 496.350000 658.500000 497.650000 ;
      RECT 616.500000 496.350000 649.500000 497.650000 ;
      RECT 607.500000 496.350000 608.500000 497.650000 ;
      RECT 566.500000 496.350000 599.500000 497.650000 ;
      RECT 557.500000 496.350000 558.500000 497.650000 ;
      RECT 516.500000 496.350000 549.500000 497.650000 ;
      RECT 507.500000 496.350000 508.500000 497.650000 ;
      RECT 466.500000 496.350000 499.500000 497.650000 ;
      RECT 457.500000 496.350000 458.500000 497.650000 ;
      RECT 416.500000 496.350000 449.500000 497.650000 ;
      RECT 407.500000 496.350000 408.500000 497.650000 ;
      RECT 396.500000 496.350000 399.500000 499.650000 ;
      RECT 382.500000 496.350000 383.500000 497.650000 ;
      RECT 357.500000 496.350000 358.500000 497.650000 ;
      RECT 316.500000 496.350000 349.500000 497.650000 ;
      RECT 307.500000 496.350000 308.500000 497.650000 ;
      RECT 266.500000 496.350000 299.500000 497.650000 ;
      RECT 257.500000 496.350000 258.500000 497.650000 ;
      RECT 216.500000 496.350000 249.500000 497.650000 ;
      RECT 207.500000 496.350000 208.500000 497.650000 ;
      RECT 166.500000 496.350000 199.500000 497.650000 ;
      RECT 157.500000 496.350000 158.500000 497.650000 ;
      RECT 116.500000 496.350000 149.500000 497.650000 ;
      RECT 107.500000 496.350000 108.500000 497.650000 ;
      RECT 66.500000 496.350000 99.500000 497.650000 ;
      RECT 57.500000 496.350000 58.500000 497.650000 ;
      RECT 29.500000 496.350000 49.500000 497.650000 ;
      RECT 15.500000 496.350000 16.500000 497.650000 ;
      RECT 0.000000 496.350000 2.500000 499.650000 ;
      RECT 1139.000000 495.650000 1158.500000 496.350000 ;
      RECT 716.500000 495.650000 749.000000 496.350000 ;
      RECT 666.500000 495.650000 708.500000 496.350000 ;
      RECT 616.500000 495.650000 658.500000 496.350000 ;
      RECT 566.500000 495.650000 608.500000 496.350000 ;
      RECT 516.500000 495.650000 558.500000 496.350000 ;
      RECT 466.500000 495.650000 508.500000 496.350000 ;
      RECT 416.500000 495.650000 458.500000 496.350000 ;
      RECT 382.500000 495.650000 408.500000 496.350000 ;
      RECT 316.500000 495.650000 358.500000 496.350000 ;
      RECT 266.500000 495.650000 308.500000 496.350000 ;
      RECT 216.500000 495.650000 258.500000 496.350000 ;
      RECT 166.500000 495.650000 208.500000 496.350000 ;
      RECT 116.500000 495.650000 158.500000 496.350000 ;
      RECT 66.500000 495.650000 108.500000 496.350000 ;
      RECT 29.500000 495.650000 58.500000 496.350000 ;
      RECT 0.000000 495.650000 16.500000 496.350000 ;
      RECT 1166.500000 494.350000 1186.000000 497.650000 ;
      RECT 1157.500000 494.350000 1158.500000 495.650000 ;
      RECT 716.500000 494.350000 733.500000 495.650000 ;
      RECT 707.500000 494.350000 708.500000 495.650000 ;
      RECT 666.500000 494.350000 699.500000 495.650000 ;
      RECT 657.500000 494.350000 658.500000 495.650000 ;
      RECT 616.500000 494.350000 649.500000 495.650000 ;
      RECT 607.500000 494.350000 608.500000 495.650000 ;
      RECT 566.500000 494.350000 599.500000 495.650000 ;
      RECT 557.500000 494.350000 558.500000 495.650000 ;
      RECT 516.500000 494.350000 549.500000 495.650000 ;
      RECT 507.500000 494.350000 508.500000 495.650000 ;
      RECT 466.500000 494.350000 499.500000 495.650000 ;
      RECT 457.500000 494.350000 458.500000 495.650000 ;
      RECT 416.500000 494.350000 449.500000 495.650000 ;
      RECT 407.500000 494.350000 408.500000 495.650000 ;
      RECT 382.500000 494.350000 383.500000 495.650000 ;
      RECT 366.500000 494.350000 369.500000 497.650000 ;
      RECT 357.500000 494.350000 358.500000 495.650000 ;
      RECT 316.500000 494.350000 349.500000 495.650000 ;
      RECT 307.500000 494.350000 308.500000 495.650000 ;
      RECT 266.500000 494.350000 299.500000 495.650000 ;
      RECT 257.500000 494.350000 258.500000 495.650000 ;
      RECT 216.500000 494.350000 249.500000 495.650000 ;
      RECT 207.500000 494.350000 208.500000 495.650000 ;
      RECT 166.500000 494.350000 199.500000 495.650000 ;
      RECT 157.500000 494.350000 158.500000 495.650000 ;
      RECT 116.500000 494.350000 149.500000 495.650000 ;
      RECT 107.500000 494.350000 108.500000 495.650000 ;
      RECT 66.500000 494.350000 99.500000 495.650000 ;
      RECT 57.500000 494.350000 58.500000 495.650000 ;
      RECT 29.500000 494.350000 49.500000 495.650000 ;
      RECT 15.500000 494.350000 16.500000 495.650000 ;
      RECT 1157.500000 493.650000 1186.000000 494.350000 ;
      RECT 707.500000 493.650000 733.500000 494.350000 ;
      RECT 657.500000 493.650000 699.500000 494.350000 ;
      RECT 607.500000 493.650000 649.500000 494.350000 ;
      RECT 557.500000 493.650000 599.500000 494.350000 ;
      RECT 507.500000 493.650000 549.500000 494.350000 ;
      RECT 457.500000 493.650000 499.500000 494.350000 ;
      RECT 407.500000 493.650000 449.500000 494.350000 ;
      RECT 357.500000 493.650000 383.500000 494.350000 ;
      RECT 307.500000 493.650000 349.500000 494.350000 ;
      RECT 257.500000 493.650000 299.500000 494.350000 ;
      RECT 207.500000 493.650000 249.500000 494.350000 ;
      RECT 157.500000 493.650000 199.500000 494.350000 ;
      RECT 107.500000 493.650000 149.500000 494.350000 ;
      RECT 57.500000 493.650000 99.500000 494.350000 ;
      RECT 15.500000 493.650000 49.500000 494.350000 ;
      RECT 1157.500000 492.350000 1158.500000 493.650000 ;
      RECT 1139.000000 492.350000 1149.500000 495.650000 ;
      RECT 746.500000 492.350000 749.000000 495.650000 ;
      RECT 716.500000 492.350000 733.500000 493.650000 ;
      RECT 707.500000 492.350000 708.500000 493.650000 ;
      RECT 666.500000 492.350000 699.500000 493.650000 ;
      RECT 657.500000 492.350000 658.500000 493.650000 ;
      RECT 616.500000 492.350000 649.500000 493.650000 ;
      RECT 607.500000 492.350000 608.500000 493.650000 ;
      RECT 566.500000 492.350000 599.500000 493.650000 ;
      RECT 557.500000 492.350000 558.500000 493.650000 ;
      RECT 516.500000 492.350000 549.500000 493.650000 ;
      RECT 507.500000 492.350000 508.500000 493.650000 ;
      RECT 466.500000 492.350000 499.500000 493.650000 ;
      RECT 457.500000 492.350000 458.500000 493.650000 ;
      RECT 416.500000 492.350000 449.500000 493.650000 ;
      RECT 407.500000 492.350000 408.500000 493.650000 ;
      RECT 396.500000 492.350000 399.500000 495.650000 ;
      RECT 382.500000 492.350000 383.500000 493.650000 ;
      RECT 357.500000 492.350000 358.500000 493.650000 ;
      RECT 316.500000 492.350000 349.500000 493.650000 ;
      RECT 307.500000 492.350000 308.500000 493.650000 ;
      RECT 266.500000 492.350000 299.500000 493.650000 ;
      RECT 257.500000 492.350000 258.500000 493.650000 ;
      RECT 216.500000 492.350000 249.500000 493.650000 ;
      RECT 207.500000 492.350000 208.500000 493.650000 ;
      RECT 166.500000 492.350000 199.500000 493.650000 ;
      RECT 157.500000 492.350000 158.500000 493.650000 ;
      RECT 116.500000 492.350000 149.500000 493.650000 ;
      RECT 107.500000 492.350000 108.500000 493.650000 ;
      RECT 66.500000 492.350000 99.500000 493.650000 ;
      RECT 57.500000 492.350000 58.500000 493.650000 ;
      RECT 29.500000 492.350000 49.500000 493.650000 ;
      RECT 15.500000 492.350000 16.500000 493.650000 ;
      RECT 0.000000 492.350000 2.500000 495.650000 ;
      RECT 1139.000000 491.650000 1158.500000 492.350000 ;
      RECT 716.500000 491.650000 749.000000 492.350000 ;
      RECT 666.500000 491.650000 708.500000 492.350000 ;
      RECT 616.500000 491.650000 658.500000 492.350000 ;
      RECT 566.500000 491.650000 608.500000 492.350000 ;
      RECT 516.500000 491.650000 558.500000 492.350000 ;
      RECT 466.500000 491.650000 508.500000 492.350000 ;
      RECT 416.500000 491.650000 458.500000 492.350000 ;
      RECT 382.500000 491.650000 408.500000 492.350000 ;
      RECT 316.500000 491.650000 358.500000 492.350000 ;
      RECT 266.500000 491.650000 308.500000 492.350000 ;
      RECT 216.500000 491.650000 258.500000 492.350000 ;
      RECT 166.500000 491.650000 208.500000 492.350000 ;
      RECT 116.500000 491.650000 158.500000 492.350000 ;
      RECT 66.500000 491.650000 108.500000 492.350000 ;
      RECT 29.500000 491.650000 58.500000 492.350000 ;
      RECT 0.000000 491.650000 16.500000 492.350000 ;
      RECT 1166.500000 490.350000 1186.000000 493.650000 ;
      RECT 1157.500000 490.350000 1158.500000 491.650000 ;
      RECT 716.500000 490.350000 733.500000 491.650000 ;
      RECT 707.500000 490.350000 708.500000 491.650000 ;
      RECT 666.500000 490.350000 699.500000 491.650000 ;
      RECT 657.500000 490.350000 658.500000 491.650000 ;
      RECT 616.500000 490.350000 649.500000 491.650000 ;
      RECT 607.500000 490.350000 608.500000 491.650000 ;
      RECT 566.500000 490.350000 599.500000 491.650000 ;
      RECT 557.500000 490.350000 558.500000 491.650000 ;
      RECT 516.500000 490.350000 549.500000 491.650000 ;
      RECT 507.500000 490.350000 508.500000 491.650000 ;
      RECT 466.500000 490.350000 499.500000 491.650000 ;
      RECT 457.500000 490.350000 458.500000 491.650000 ;
      RECT 416.500000 490.350000 449.500000 491.650000 ;
      RECT 407.500000 490.350000 408.500000 491.650000 ;
      RECT 382.500000 490.350000 399.500000 491.650000 ;
      RECT 366.500000 490.350000 369.500000 493.650000 ;
      RECT 357.500000 490.350000 358.500000 491.650000 ;
      RECT 316.500000 490.350000 349.500000 491.650000 ;
      RECT 307.500000 490.350000 308.500000 491.650000 ;
      RECT 266.500000 490.350000 299.500000 491.650000 ;
      RECT 257.500000 490.350000 258.500000 491.650000 ;
      RECT 216.500000 490.350000 249.500000 491.650000 ;
      RECT 207.500000 490.350000 208.500000 491.650000 ;
      RECT 166.500000 490.350000 199.500000 491.650000 ;
      RECT 157.500000 490.350000 158.500000 491.650000 ;
      RECT 116.500000 490.350000 149.500000 491.650000 ;
      RECT 107.500000 490.350000 108.500000 491.650000 ;
      RECT 66.500000 490.350000 99.500000 491.650000 ;
      RECT 57.500000 490.350000 58.500000 491.650000 ;
      RECT 29.500000 490.350000 49.500000 491.650000 ;
      RECT 15.500000 490.350000 16.500000 491.650000 ;
      RECT 1157.500000 489.650000 1186.000000 490.350000 ;
      RECT 707.500000 489.650000 733.500000 490.350000 ;
      RECT 657.500000 489.650000 699.500000 490.350000 ;
      RECT 607.500000 489.650000 649.500000 490.350000 ;
      RECT 557.500000 489.650000 599.500000 490.350000 ;
      RECT 507.500000 489.650000 549.500000 490.350000 ;
      RECT 457.500000 489.650000 499.500000 490.350000 ;
      RECT 407.500000 489.650000 449.500000 490.350000 ;
      RECT 357.500000 489.650000 399.500000 490.350000 ;
      RECT 307.500000 489.650000 349.500000 490.350000 ;
      RECT 257.500000 489.650000 299.500000 490.350000 ;
      RECT 207.500000 489.650000 249.500000 490.350000 ;
      RECT 157.500000 489.650000 199.500000 490.350000 ;
      RECT 107.500000 489.650000 149.500000 490.350000 ;
      RECT 57.500000 489.650000 99.500000 490.350000 ;
      RECT 15.500000 489.650000 49.500000 490.350000 ;
      RECT 1157.500000 488.350000 1158.500000 489.650000 ;
      RECT 1139.000000 488.350000 1149.500000 491.650000 ;
      RECT 746.500000 488.350000 749.000000 491.650000 ;
      RECT 732.500000 488.350000 733.500000 489.650000 ;
      RECT 707.500000 488.350000 708.500000 489.650000 ;
      RECT 666.500000 488.350000 699.500000 489.650000 ;
      RECT 657.500000 488.350000 658.500000 489.650000 ;
      RECT 616.500000 488.350000 649.500000 489.650000 ;
      RECT 607.500000 488.350000 608.500000 489.650000 ;
      RECT 566.500000 488.350000 599.500000 489.650000 ;
      RECT 557.500000 488.350000 558.500000 489.650000 ;
      RECT 516.500000 488.350000 549.500000 489.650000 ;
      RECT 507.500000 488.350000 508.500000 489.650000 ;
      RECT 466.500000 488.350000 499.500000 489.650000 ;
      RECT 457.500000 488.350000 458.500000 489.650000 ;
      RECT 416.500000 488.350000 449.500000 489.650000 ;
      RECT 407.500000 488.350000 408.500000 489.650000 ;
      RECT 382.500000 488.350000 399.500000 489.650000 ;
      RECT 357.500000 488.350000 358.500000 489.650000 ;
      RECT 316.500000 488.350000 349.500000 489.650000 ;
      RECT 307.500000 488.350000 308.500000 489.650000 ;
      RECT 266.500000 488.350000 299.500000 489.650000 ;
      RECT 257.500000 488.350000 258.500000 489.650000 ;
      RECT 216.500000 488.350000 249.500000 489.650000 ;
      RECT 207.500000 488.350000 208.500000 489.650000 ;
      RECT 166.500000 488.350000 199.500000 489.650000 ;
      RECT 157.500000 488.350000 158.500000 489.650000 ;
      RECT 116.500000 488.350000 149.500000 489.650000 ;
      RECT 107.500000 488.350000 108.500000 489.650000 ;
      RECT 66.500000 488.350000 99.500000 489.650000 ;
      RECT 57.500000 488.350000 58.500000 489.650000 ;
      RECT 29.500000 488.350000 49.500000 489.650000 ;
      RECT 15.500000 488.350000 16.500000 489.650000 ;
      RECT 0.000000 488.350000 2.500000 491.650000 ;
      RECT 1139.000000 487.650000 1158.500000 488.350000 ;
      RECT 732.500000 487.650000 749.000000 488.350000 ;
      RECT 666.500000 487.650000 708.500000 488.350000 ;
      RECT 616.500000 487.650000 658.500000 488.350000 ;
      RECT 566.500000 487.650000 608.500000 488.350000 ;
      RECT 516.500000 487.650000 558.500000 488.350000 ;
      RECT 466.500000 487.650000 508.500000 488.350000 ;
      RECT 416.500000 487.650000 458.500000 488.350000 ;
      RECT 382.500000 487.650000 408.500000 488.350000 ;
      RECT 316.500000 487.650000 358.500000 488.350000 ;
      RECT 266.500000 487.650000 308.500000 488.350000 ;
      RECT 216.500000 487.650000 258.500000 488.350000 ;
      RECT 166.500000 487.650000 208.500000 488.350000 ;
      RECT 116.500000 487.650000 158.500000 488.350000 ;
      RECT 66.500000 487.650000 108.500000 488.350000 ;
      RECT 29.500000 487.650000 58.500000 488.350000 ;
      RECT 0.000000 487.650000 16.500000 488.350000 ;
      RECT 1166.500000 486.350000 1186.000000 489.650000 ;
      RECT 1157.500000 486.350000 1158.500000 487.650000 ;
      RECT 732.500000 486.350000 733.500000 487.650000 ;
      RECT 716.500000 486.350000 719.500000 489.650000 ;
      RECT 707.500000 486.350000 708.500000 487.650000 ;
      RECT 666.500000 486.350000 699.500000 487.650000 ;
      RECT 657.500000 486.350000 658.500000 487.650000 ;
      RECT 616.500000 486.350000 649.500000 487.650000 ;
      RECT 607.500000 486.350000 608.500000 487.650000 ;
      RECT 566.500000 486.350000 599.500000 487.650000 ;
      RECT 557.500000 486.350000 558.500000 487.650000 ;
      RECT 516.500000 486.350000 549.500000 487.650000 ;
      RECT 507.500000 486.350000 508.500000 487.650000 ;
      RECT 466.500000 486.350000 499.500000 487.650000 ;
      RECT 457.500000 486.350000 458.500000 487.650000 ;
      RECT 416.500000 486.350000 449.500000 487.650000 ;
      RECT 407.500000 486.350000 408.500000 487.650000 ;
      RECT 382.500000 486.350000 399.500000 487.650000 ;
      RECT 366.500000 486.350000 369.500000 489.650000 ;
      RECT 357.500000 486.350000 358.500000 487.650000 ;
      RECT 316.500000 486.350000 349.500000 487.650000 ;
      RECT 307.500000 486.350000 308.500000 487.650000 ;
      RECT 266.500000 486.350000 299.500000 487.650000 ;
      RECT 257.500000 486.350000 258.500000 487.650000 ;
      RECT 216.500000 486.350000 249.500000 487.650000 ;
      RECT 207.500000 486.350000 208.500000 487.650000 ;
      RECT 166.500000 486.350000 199.500000 487.650000 ;
      RECT 157.500000 486.350000 158.500000 487.650000 ;
      RECT 116.500000 486.350000 149.500000 487.650000 ;
      RECT 107.500000 486.350000 108.500000 487.650000 ;
      RECT 66.500000 486.350000 99.500000 487.650000 ;
      RECT 57.500000 486.350000 58.500000 487.650000 ;
      RECT 29.500000 486.350000 49.500000 487.650000 ;
      RECT 15.500000 486.350000 16.500000 487.650000 ;
      RECT 1157.500000 485.650000 1186.000000 486.350000 ;
      RECT 707.500000 485.650000 733.500000 486.350000 ;
      RECT 657.500000 485.650000 699.500000 486.350000 ;
      RECT 607.500000 485.650000 649.500000 486.350000 ;
      RECT 557.500000 485.650000 599.500000 486.350000 ;
      RECT 507.500000 485.650000 549.500000 486.350000 ;
      RECT 457.500000 485.650000 499.500000 486.350000 ;
      RECT 407.500000 485.650000 449.500000 486.350000 ;
      RECT 357.500000 485.650000 399.500000 486.350000 ;
      RECT 307.500000 485.650000 349.500000 486.350000 ;
      RECT 257.500000 485.650000 299.500000 486.350000 ;
      RECT 207.500000 485.650000 249.500000 486.350000 ;
      RECT 157.500000 485.650000 199.500000 486.350000 ;
      RECT 107.500000 485.650000 149.500000 486.350000 ;
      RECT 57.500000 485.650000 99.500000 486.350000 ;
      RECT 15.500000 485.650000 49.500000 486.350000 ;
      RECT 1157.500000 484.350000 1158.500000 485.650000 ;
      RECT 1139.000000 484.350000 1149.500000 487.650000 ;
      RECT 746.500000 484.350000 749.000000 487.650000 ;
      RECT 732.500000 484.350000 733.500000 485.650000 ;
      RECT 707.500000 484.350000 708.500000 485.650000 ;
      RECT 666.500000 484.350000 699.500000 485.650000 ;
      RECT 657.500000 484.350000 658.500000 485.650000 ;
      RECT 616.500000 484.350000 649.500000 485.650000 ;
      RECT 607.500000 484.350000 608.500000 485.650000 ;
      RECT 566.500000 484.350000 599.500000 485.650000 ;
      RECT 557.500000 484.350000 558.500000 485.650000 ;
      RECT 516.500000 484.350000 549.500000 485.650000 ;
      RECT 507.500000 484.350000 508.500000 485.650000 ;
      RECT 466.500000 484.350000 499.500000 485.650000 ;
      RECT 457.500000 484.350000 458.500000 485.650000 ;
      RECT 416.500000 484.350000 449.500000 485.650000 ;
      RECT 407.500000 484.350000 408.500000 485.650000 ;
      RECT 382.500000 484.350000 399.500000 485.650000 ;
      RECT 357.500000 484.350000 358.500000 485.650000 ;
      RECT 316.500000 484.350000 349.500000 485.650000 ;
      RECT 307.500000 484.350000 308.500000 485.650000 ;
      RECT 266.500000 484.350000 299.500000 485.650000 ;
      RECT 257.500000 484.350000 258.500000 485.650000 ;
      RECT 216.500000 484.350000 249.500000 485.650000 ;
      RECT 207.500000 484.350000 208.500000 485.650000 ;
      RECT 166.500000 484.350000 199.500000 485.650000 ;
      RECT 157.500000 484.350000 158.500000 485.650000 ;
      RECT 116.500000 484.350000 149.500000 485.650000 ;
      RECT 107.500000 484.350000 108.500000 485.650000 ;
      RECT 66.500000 484.350000 99.500000 485.650000 ;
      RECT 57.500000 484.350000 58.500000 485.650000 ;
      RECT 29.500000 484.350000 49.500000 485.650000 ;
      RECT 15.500000 484.350000 16.500000 485.650000 ;
      RECT 0.000000 484.350000 2.500000 487.650000 ;
      RECT 1139.000000 483.650000 1158.500000 484.350000 ;
      RECT 732.500000 483.650000 749.000000 484.350000 ;
      RECT 666.500000 483.650000 708.500000 484.350000 ;
      RECT 616.500000 483.650000 658.500000 484.350000 ;
      RECT 566.500000 483.650000 608.500000 484.350000 ;
      RECT 516.500000 483.650000 558.500000 484.350000 ;
      RECT 466.500000 483.650000 508.500000 484.350000 ;
      RECT 416.500000 483.650000 458.500000 484.350000 ;
      RECT 382.500000 483.650000 408.500000 484.350000 ;
      RECT 316.500000 483.650000 358.500000 484.350000 ;
      RECT 266.500000 483.650000 308.500000 484.350000 ;
      RECT 216.500000 483.650000 258.500000 484.350000 ;
      RECT 166.500000 483.650000 208.500000 484.350000 ;
      RECT 116.500000 483.650000 158.500000 484.350000 ;
      RECT 66.500000 483.650000 108.500000 484.350000 ;
      RECT 29.500000 483.650000 58.500000 484.350000 ;
      RECT 0.000000 483.650000 16.500000 484.350000 ;
      RECT 1166.500000 482.350000 1186.000000 485.650000 ;
      RECT 1157.500000 482.350000 1158.500000 483.650000 ;
      RECT 732.500000 482.350000 733.500000 483.650000 ;
      RECT 716.500000 482.350000 719.500000 485.650000 ;
      RECT 707.500000 482.350000 708.500000 483.650000 ;
      RECT 666.500000 482.350000 699.500000 483.650000 ;
      RECT 657.500000 482.350000 658.500000 483.650000 ;
      RECT 616.500000 482.350000 649.500000 483.650000 ;
      RECT 607.500000 482.350000 608.500000 483.650000 ;
      RECT 566.500000 482.350000 599.500000 483.650000 ;
      RECT 557.500000 482.350000 558.500000 483.650000 ;
      RECT 516.500000 482.350000 549.500000 483.650000 ;
      RECT 507.500000 482.350000 508.500000 483.650000 ;
      RECT 466.500000 482.350000 499.500000 483.650000 ;
      RECT 457.500000 482.350000 458.500000 483.650000 ;
      RECT 416.500000 482.350000 449.500000 483.650000 ;
      RECT 407.500000 482.350000 408.500000 483.650000 ;
      RECT 382.500000 482.350000 399.500000 483.650000 ;
      RECT 366.500000 482.350000 369.500000 485.650000 ;
      RECT 357.500000 482.350000 358.500000 483.650000 ;
      RECT 316.500000 482.350000 349.500000 483.650000 ;
      RECT 307.500000 482.350000 308.500000 483.650000 ;
      RECT 266.500000 482.350000 299.500000 483.650000 ;
      RECT 257.500000 482.350000 258.500000 483.650000 ;
      RECT 216.500000 482.350000 249.500000 483.650000 ;
      RECT 207.500000 482.350000 208.500000 483.650000 ;
      RECT 166.500000 482.350000 199.500000 483.650000 ;
      RECT 157.500000 482.350000 158.500000 483.650000 ;
      RECT 116.500000 482.350000 149.500000 483.650000 ;
      RECT 107.500000 482.350000 108.500000 483.650000 ;
      RECT 66.500000 482.350000 99.500000 483.650000 ;
      RECT 57.500000 482.350000 58.500000 483.650000 ;
      RECT 29.500000 482.350000 49.500000 483.650000 ;
      RECT 15.500000 482.350000 16.500000 483.650000 ;
      RECT 1157.500000 481.650000 1186.000000 482.350000 ;
      RECT 707.500000 481.650000 733.500000 482.350000 ;
      RECT 657.500000 481.650000 699.500000 482.350000 ;
      RECT 607.500000 481.650000 649.500000 482.350000 ;
      RECT 557.500000 481.650000 599.500000 482.350000 ;
      RECT 507.500000 481.650000 549.500000 482.350000 ;
      RECT 457.500000 481.650000 499.500000 482.350000 ;
      RECT 407.500000 481.650000 449.500000 482.350000 ;
      RECT 357.500000 481.650000 399.500000 482.350000 ;
      RECT 307.500000 481.650000 349.500000 482.350000 ;
      RECT 257.500000 481.650000 299.500000 482.350000 ;
      RECT 207.500000 481.650000 249.500000 482.350000 ;
      RECT 157.500000 481.650000 199.500000 482.350000 ;
      RECT 107.500000 481.650000 149.500000 482.350000 ;
      RECT 57.500000 481.650000 99.500000 482.350000 ;
      RECT 15.500000 481.650000 49.500000 482.350000 ;
      RECT 1157.500000 480.350000 1158.500000 481.650000 ;
      RECT 1139.000000 480.350000 1149.500000 483.650000 ;
      RECT 746.500000 480.350000 749.000000 483.650000 ;
      RECT 732.500000 480.350000 733.500000 481.650000 ;
      RECT 707.500000 480.350000 708.500000 481.650000 ;
      RECT 666.500000 480.350000 699.500000 481.650000 ;
      RECT 657.500000 480.350000 658.500000 481.650000 ;
      RECT 616.500000 480.350000 649.500000 481.650000 ;
      RECT 607.500000 480.350000 608.500000 481.650000 ;
      RECT 566.500000 480.350000 599.500000 481.650000 ;
      RECT 557.500000 480.350000 558.500000 481.650000 ;
      RECT 516.500000 480.350000 549.500000 481.650000 ;
      RECT 507.500000 480.350000 508.500000 481.650000 ;
      RECT 466.500000 480.350000 499.500000 481.650000 ;
      RECT 457.500000 480.350000 458.500000 481.650000 ;
      RECT 416.500000 480.350000 449.500000 481.650000 ;
      RECT 407.500000 480.350000 408.500000 481.650000 ;
      RECT 382.500000 480.350000 399.500000 481.650000 ;
      RECT 357.500000 480.350000 358.500000 481.650000 ;
      RECT 316.500000 480.350000 349.500000 481.650000 ;
      RECT 307.500000 480.350000 308.500000 481.650000 ;
      RECT 266.500000 480.350000 299.500000 481.650000 ;
      RECT 257.500000 480.350000 258.500000 481.650000 ;
      RECT 216.500000 480.350000 249.500000 481.650000 ;
      RECT 207.500000 480.350000 208.500000 481.650000 ;
      RECT 166.500000 480.350000 199.500000 481.650000 ;
      RECT 157.500000 480.350000 158.500000 481.650000 ;
      RECT 116.500000 480.350000 149.500000 481.650000 ;
      RECT 107.500000 480.350000 108.500000 481.650000 ;
      RECT 66.500000 480.350000 99.500000 481.650000 ;
      RECT 57.500000 480.350000 58.500000 481.650000 ;
      RECT 29.500000 480.350000 49.500000 481.650000 ;
      RECT 15.500000 480.350000 16.500000 481.650000 ;
      RECT 0.000000 480.350000 2.500000 483.650000 ;
      RECT 1139.000000 479.650000 1158.500000 480.350000 ;
      RECT 732.500000 479.650000 749.000000 480.350000 ;
      RECT 666.500000 479.650000 708.500000 480.350000 ;
      RECT 616.500000 479.650000 658.500000 480.350000 ;
      RECT 566.500000 479.650000 608.500000 480.350000 ;
      RECT 516.500000 479.650000 558.500000 480.350000 ;
      RECT 466.500000 479.650000 508.500000 480.350000 ;
      RECT 416.500000 479.650000 458.500000 480.350000 ;
      RECT 382.500000 479.650000 408.500000 480.350000 ;
      RECT 316.500000 479.650000 358.500000 480.350000 ;
      RECT 266.500000 479.650000 308.500000 480.350000 ;
      RECT 216.500000 479.650000 258.500000 480.350000 ;
      RECT 166.500000 479.650000 208.500000 480.350000 ;
      RECT 116.500000 479.650000 158.500000 480.350000 ;
      RECT 66.500000 479.650000 108.500000 480.350000 ;
      RECT 29.500000 479.650000 58.500000 480.350000 ;
      RECT 0.000000 479.650000 16.500000 480.350000 ;
      RECT 1166.500000 478.350000 1186.000000 481.650000 ;
      RECT 1157.500000 478.350000 1158.500000 479.650000 ;
      RECT 732.500000 478.350000 733.500000 479.650000 ;
      RECT 716.500000 478.350000 719.500000 481.650000 ;
      RECT 707.500000 478.350000 708.500000 479.650000 ;
      RECT 666.500000 478.350000 699.500000 479.650000 ;
      RECT 657.500000 478.350000 658.500000 479.650000 ;
      RECT 616.500000 478.350000 649.500000 479.650000 ;
      RECT 607.500000 478.350000 608.500000 479.650000 ;
      RECT 566.500000 478.350000 599.500000 479.650000 ;
      RECT 557.500000 478.350000 558.500000 479.650000 ;
      RECT 516.500000 478.350000 549.500000 479.650000 ;
      RECT 507.500000 478.350000 508.500000 479.650000 ;
      RECT 466.500000 478.350000 499.500000 479.650000 ;
      RECT 457.500000 478.350000 458.500000 479.650000 ;
      RECT 416.500000 478.350000 449.500000 479.650000 ;
      RECT 407.500000 478.350000 408.500000 479.650000 ;
      RECT 382.500000 478.350000 399.500000 479.650000 ;
      RECT 366.500000 478.350000 369.500000 481.650000 ;
      RECT 357.500000 478.350000 358.500000 479.650000 ;
      RECT 316.500000 478.350000 349.500000 479.650000 ;
      RECT 307.500000 478.350000 308.500000 479.650000 ;
      RECT 266.500000 478.350000 299.500000 479.650000 ;
      RECT 257.500000 478.350000 258.500000 479.650000 ;
      RECT 216.500000 478.350000 249.500000 479.650000 ;
      RECT 207.500000 478.350000 208.500000 479.650000 ;
      RECT 166.500000 478.350000 199.500000 479.650000 ;
      RECT 157.500000 478.350000 158.500000 479.650000 ;
      RECT 116.500000 478.350000 149.500000 479.650000 ;
      RECT 107.500000 478.350000 108.500000 479.650000 ;
      RECT 66.500000 478.350000 99.500000 479.650000 ;
      RECT 57.500000 478.350000 58.500000 479.650000 ;
      RECT 29.500000 478.350000 49.500000 479.650000 ;
      RECT 15.500000 478.350000 16.500000 479.650000 ;
      RECT 1157.500000 477.650000 1186.000000 478.350000 ;
      RECT 707.500000 477.650000 733.500000 478.350000 ;
      RECT 657.500000 477.650000 699.500000 478.350000 ;
      RECT 607.500000 477.650000 649.500000 478.350000 ;
      RECT 557.500000 477.650000 599.500000 478.350000 ;
      RECT 507.500000 477.650000 549.500000 478.350000 ;
      RECT 457.500000 477.650000 499.500000 478.350000 ;
      RECT 407.500000 477.650000 449.500000 478.350000 ;
      RECT 357.500000 477.650000 399.500000 478.350000 ;
      RECT 307.500000 477.650000 349.500000 478.350000 ;
      RECT 257.500000 477.650000 299.500000 478.350000 ;
      RECT 207.500000 477.650000 249.500000 478.350000 ;
      RECT 157.500000 477.650000 199.500000 478.350000 ;
      RECT 107.500000 477.650000 149.500000 478.350000 ;
      RECT 57.500000 477.650000 99.500000 478.350000 ;
      RECT 15.500000 477.650000 49.500000 478.350000 ;
      RECT 1157.500000 476.350000 1158.500000 477.650000 ;
      RECT 1139.000000 476.350000 1149.500000 479.650000 ;
      RECT 746.500000 476.350000 749.000000 479.650000 ;
      RECT 732.500000 476.350000 733.500000 477.650000 ;
      RECT 707.500000 476.350000 708.500000 477.650000 ;
      RECT 666.500000 476.350000 699.500000 477.650000 ;
      RECT 657.500000 476.350000 658.500000 477.650000 ;
      RECT 616.500000 476.350000 649.500000 477.650000 ;
      RECT 607.500000 476.350000 608.500000 477.650000 ;
      RECT 566.500000 476.350000 599.500000 477.650000 ;
      RECT 557.500000 476.350000 558.500000 477.650000 ;
      RECT 516.500000 476.350000 549.500000 477.650000 ;
      RECT 507.500000 476.350000 508.500000 477.650000 ;
      RECT 466.500000 476.350000 499.500000 477.650000 ;
      RECT 457.500000 476.350000 458.500000 477.650000 ;
      RECT 416.500000 476.350000 449.500000 477.650000 ;
      RECT 407.500000 476.350000 408.500000 477.650000 ;
      RECT 366.500000 476.350000 399.500000 477.650000 ;
      RECT 357.500000 476.350000 358.500000 477.650000 ;
      RECT 316.500000 476.350000 349.500000 477.650000 ;
      RECT 307.500000 476.350000 308.500000 477.650000 ;
      RECT 266.500000 476.350000 299.500000 477.650000 ;
      RECT 257.500000 476.350000 258.500000 477.650000 ;
      RECT 216.500000 476.350000 249.500000 477.650000 ;
      RECT 207.500000 476.350000 208.500000 477.650000 ;
      RECT 166.500000 476.350000 199.500000 477.650000 ;
      RECT 157.500000 476.350000 158.500000 477.650000 ;
      RECT 116.500000 476.350000 149.500000 477.650000 ;
      RECT 107.500000 476.350000 108.500000 477.650000 ;
      RECT 66.500000 476.350000 99.500000 477.650000 ;
      RECT 57.500000 476.350000 58.500000 477.650000 ;
      RECT 29.500000 476.350000 49.500000 477.650000 ;
      RECT 15.500000 476.350000 16.500000 477.650000 ;
      RECT 0.000000 476.350000 2.500000 479.650000 ;
      RECT 1139.000000 475.650000 1158.500000 476.350000 ;
      RECT 732.500000 475.650000 749.000000 476.350000 ;
      RECT 666.500000 475.650000 708.500000 476.350000 ;
      RECT 616.500000 475.650000 658.500000 476.350000 ;
      RECT 566.500000 475.650000 608.500000 476.350000 ;
      RECT 516.500000 475.650000 558.500000 476.350000 ;
      RECT 466.500000 475.650000 508.500000 476.350000 ;
      RECT 416.500000 475.650000 458.500000 476.350000 ;
      RECT 366.500000 475.650000 408.500000 476.350000 ;
      RECT 316.500000 475.650000 358.500000 476.350000 ;
      RECT 266.500000 475.650000 308.500000 476.350000 ;
      RECT 216.500000 475.650000 258.500000 476.350000 ;
      RECT 166.500000 475.650000 208.500000 476.350000 ;
      RECT 116.500000 475.650000 158.500000 476.350000 ;
      RECT 66.500000 475.650000 108.500000 476.350000 ;
      RECT 29.500000 475.650000 58.500000 476.350000 ;
      RECT 0.000000 475.650000 16.500000 476.350000 ;
      RECT 1166.500000 474.350000 1186.000000 477.650000 ;
      RECT 1157.500000 474.350000 1158.500000 475.650000 ;
      RECT 732.500000 474.350000 733.500000 475.650000 ;
      RECT 716.500000 474.350000 719.500000 477.650000 ;
      RECT 707.500000 474.350000 708.500000 475.650000 ;
      RECT 666.500000 474.350000 699.500000 475.650000 ;
      RECT 657.500000 474.350000 658.500000 475.650000 ;
      RECT 616.500000 474.350000 649.500000 475.650000 ;
      RECT 607.500000 474.350000 608.500000 475.650000 ;
      RECT 566.500000 474.350000 599.500000 475.650000 ;
      RECT 557.500000 474.350000 558.500000 475.650000 ;
      RECT 516.500000 474.350000 549.500000 475.650000 ;
      RECT 507.500000 474.350000 508.500000 475.650000 ;
      RECT 466.500000 474.350000 499.500000 475.650000 ;
      RECT 457.500000 474.350000 458.500000 475.650000 ;
      RECT 416.500000 474.350000 449.500000 475.650000 ;
      RECT 407.500000 474.350000 408.500000 475.650000 ;
      RECT 366.500000 474.350000 399.500000 475.650000 ;
      RECT 357.500000 474.350000 358.500000 475.650000 ;
      RECT 316.500000 474.350000 349.500000 475.650000 ;
      RECT 307.500000 474.350000 308.500000 475.650000 ;
      RECT 266.500000 474.350000 299.500000 475.650000 ;
      RECT 257.500000 474.350000 258.500000 475.650000 ;
      RECT 216.500000 474.350000 249.500000 475.650000 ;
      RECT 207.500000 474.350000 208.500000 475.650000 ;
      RECT 166.500000 474.350000 199.500000 475.650000 ;
      RECT 157.500000 474.350000 158.500000 475.650000 ;
      RECT 116.500000 474.350000 149.500000 475.650000 ;
      RECT 107.500000 474.350000 108.500000 475.650000 ;
      RECT 66.500000 474.350000 99.500000 475.650000 ;
      RECT 57.500000 474.350000 58.500000 475.650000 ;
      RECT 29.500000 474.350000 49.500000 475.650000 ;
      RECT 15.500000 474.350000 16.500000 475.650000 ;
      RECT 1157.500000 473.650000 1186.000000 474.350000 ;
      RECT 707.500000 473.650000 733.500000 474.350000 ;
      RECT 657.500000 473.650000 699.500000 474.350000 ;
      RECT 607.500000 473.650000 649.500000 474.350000 ;
      RECT 557.500000 473.650000 599.500000 474.350000 ;
      RECT 507.500000 473.650000 549.500000 474.350000 ;
      RECT 457.500000 473.650000 499.500000 474.350000 ;
      RECT 407.500000 473.650000 449.500000 474.350000 ;
      RECT 357.500000 473.650000 399.500000 474.350000 ;
      RECT 307.500000 473.650000 349.500000 474.350000 ;
      RECT 257.500000 473.650000 299.500000 474.350000 ;
      RECT 207.500000 473.650000 249.500000 474.350000 ;
      RECT 157.500000 473.650000 199.500000 474.350000 ;
      RECT 107.500000 473.650000 149.500000 474.350000 ;
      RECT 57.500000 473.650000 99.500000 474.350000 ;
      RECT 15.500000 473.650000 49.500000 474.350000 ;
      RECT 1157.500000 472.350000 1158.500000 473.650000 ;
      RECT 1139.000000 472.350000 1149.500000 475.650000 ;
      RECT 746.500000 472.350000 749.000000 475.650000 ;
      RECT 732.500000 472.350000 733.500000 473.650000 ;
      RECT 707.500000 472.350000 708.500000 473.650000 ;
      RECT 666.500000 472.350000 699.500000 473.650000 ;
      RECT 657.500000 472.350000 658.500000 473.650000 ;
      RECT 616.500000 472.350000 649.500000 473.650000 ;
      RECT 607.500000 472.350000 608.500000 473.650000 ;
      RECT 566.500000 472.350000 599.500000 473.650000 ;
      RECT 557.500000 472.350000 558.500000 473.650000 ;
      RECT 516.500000 472.350000 549.500000 473.650000 ;
      RECT 507.500000 472.350000 508.500000 473.650000 ;
      RECT 466.500000 472.350000 499.500000 473.650000 ;
      RECT 457.500000 472.350000 458.500000 473.650000 ;
      RECT 416.500000 472.350000 449.500000 473.650000 ;
      RECT 407.500000 472.350000 408.500000 473.650000 ;
      RECT 366.500000 472.350000 399.500000 473.650000 ;
      RECT 357.500000 472.350000 358.500000 473.650000 ;
      RECT 316.500000 472.350000 349.500000 473.650000 ;
      RECT 307.500000 472.350000 308.500000 473.650000 ;
      RECT 266.500000 472.350000 299.500000 473.650000 ;
      RECT 257.500000 472.350000 258.500000 473.650000 ;
      RECT 216.500000 472.350000 249.500000 473.650000 ;
      RECT 207.500000 472.350000 208.500000 473.650000 ;
      RECT 166.500000 472.350000 199.500000 473.650000 ;
      RECT 157.500000 472.350000 158.500000 473.650000 ;
      RECT 116.500000 472.350000 149.500000 473.650000 ;
      RECT 107.500000 472.350000 108.500000 473.650000 ;
      RECT 66.500000 472.350000 99.500000 473.650000 ;
      RECT 57.500000 472.350000 58.500000 473.650000 ;
      RECT 29.500000 472.350000 49.500000 473.650000 ;
      RECT 15.500000 472.350000 16.500000 473.650000 ;
      RECT 0.000000 472.350000 2.500000 475.650000 ;
      RECT 1139.000000 471.650000 1158.500000 472.350000 ;
      RECT 732.500000 471.650000 749.000000 472.350000 ;
      RECT 666.500000 471.650000 708.500000 472.350000 ;
      RECT 616.500000 471.650000 658.500000 472.350000 ;
      RECT 566.500000 471.650000 608.500000 472.350000 ;
      RECT 516.500000 471.650000 558.500000 472.350000 ;
      RECT 466.500000 471.650000 508.500000 472.350000 ;
      RECT 416.500000 471.650000 458.500000 472.350000 ;
      RECT 366.500000 471.650000 408.500000 472.350000 ;
      RECT 316.500000 471.650000 358.500000 472.350000 ;
      RECT 266.500000 471.650000 308.500000 472.350000 ;
      RECT 216.500000 471.650000 258.500000 472.350000 ;
      RECT 166.500000 471.650000 208.500000 472.350000 ;
      RECT 116.500000 471.650000 158.500000 472.350000 ;
      RECT 66.500000 471.650000 108.500000 472.350000 ;
      RECT 29.500000 471.650000 58.500000 472.350000 ;
      RECT 0.000000 471.650000 16.500000 472.350000 ;
      RECT 1166.500000 470.350000 1186.000000 473.650000 ;
      RECT 1157.500000 470.350000 1158.500000 471.650000 ;
      RECT 732.500000 470.350000 733.500000 471.650000 ;
      RECT 716.500000 470.350000 719.500000 473.650000 ;
      RECT 707.500000 470.350000 708.500000 471.650000 ;
      RECT 666.500000 470.350000 699.500000 471.650000 ;
      RECT 657.500000 470.350000 658.500000 471.650000 ;
      RECT 616.500000 470.350000 649.500000 471.650000 ;
      RECT 607.500000 470.350000 608.500000 471.650000 ;
      RECT 566.500000 470.350000 599.500000 471.650000 ;
      RECT 557.500000 470.350000 558.500000 471.650000 ;
      RECT 516.500000 470.350000 549.500000 471.650000 ;
      RECT 507.500000 470.350000 508.500000 471.650000 ;
      RECT 466.500000 470.350000 499.500000 471.650000 ;
      RECT 457.500000 470.350000 458.500000 471.650000 ;
      RECT 416.500000 470.350000 449.500000 471.650000 ;
      RECT 407.500000 470.350000 408.500000 471.650000 ;
      RECT 366.500000 470.350000 399.500000 471.650000 ;
      RECT 357.500000 470.350000 358.500000 471.650000 ;
      RECT 316.500000 470.350000 349.500000 471.650000 ;
      RECT 307.500000 470.350000 308.500000 471.650000 ;
      RECT 266.500000 470.350000 299.500000 471.650000 ;
      RECT 257.500000 470.350000 258.500000 471.650000 ;
      RECT 216.500000 470.350000 249.500000 471.650000 ;
      RECT 207.500000 470.350000 208.500000 471.650000 ;
      RECT 166.500000 470.350000 199.500000 471.650000 ;
      RECT 157.500000 470.350000 158.500000 471.650000 ;
      RECT 116.500000 470.350000 149.500000 471.650000 ;
      RECT 107.500000 470.350000 108.500000 471.650000 ;
      RECT 66.500000 470.350000 99.500000 471.650000 ;
      RECT 57.500000 470.350000 58.500000 471.650000 ;
      RECT 29.500000 470.350000 49.500000 471.650000 ;
      RECT 15.500000 470.350000 16.500000 471.650000 ;
      RECT 1157.500000 469.650000 1186.000000 470.350000 ;
      RECT 707.500000 469.650000 733.500000 470.350000 ;
      RECT 657.500000 469.650000 699.500000 470.350000 ;
      RECT 607.500000 469.650000 649.500000 470.350000 ;
      RECT 557.500000 469.650000 599.500000 470.350000 ;
      RECT 507.500000 469.650000 549.500000 470.350000 ;
      RECT 457.500000 469.650000 499.500000 470.350000 ;
      RECT 407.500000 469.650000 449.500000 470.350000 ;
      RECT 357.500000 469.650000 399.500000 470.350000 ;
      RECT 307.500000 469.650000 349.500000 470.350000 ;
      RECT 257.500000 469.650000 299.500000 470.350000 ;
      RECT 207.500000 469.650000 249.500000 470.350000 ;
      RECT 157.500000 469.650000 199.500000 470.350000 ;
      RECT 107.500000 469.650000 149.500000 470.350000 ;
      RECT 57.500000 469.650000 99.500000 470.350000 ;
      RECT 15.500000 469.650000 49.500000 470.350000 ;
      RECT 1157.500000 468.350000 1158.500000 469.650000 ;
      RECT 1139.000000 468.350000 1149.500000 471.650000 ;
      RECT 746.500000 468.350000 749.000000 471.650000 ;
      RECT 732.500000 468.350000 733.500000 469.650000 ;
      RECT 707.500000 468.350000 708.500000 469.650000 ;
      RECT 666.500000 468.350000 699.500000 469.650000 ;
      RECT 657.500000 468.350000 658.500000 469.650000 ;
      RECT 616.500000 468.350000 649.500000 469.650000 ;
      RECT 607.500000 468.350000 608.500000 469.650000 ;
      RECT 566.500000 468.350000 599.500000 469.650000 ;
      RECT 557.500000 468.350000 558.500000 469.650000 ;
      RECT 516.500000 468.350000 549.500000 469.650000 ;
      RECT 507.500000 468.350000 508.500000 469.650000 ;
      RECT 466.500000 468.350000 499.500000 469.650000 ;
      RECT 457.500000 468.350000 458.500000 469.650000 ;
      RECT 416.500000 468.350000 449.500000 469.650000 ;
      RECT 407.500000 468.350000 408.500000 469.650000 ;
      RECT 366.500000 468.350000 399.500000 469.650000 ;
      RECT 357.500000 468.350000 358.500000 469.650000 ;
      RECT 316.500000 468.350000 349.500000 469.650000 ;
      RECT 307.500000 468.350000 308.500000 469.650000 ;
      RECT 266.500000 468.350000 299.500000 469.650000 ;
      RECT 257.500000 468.350000 258.500000 469.650000 ;
      RECT 216.500000 468.350000 249.500000 469.650000 ;
      RECT 207.500000 468.350000 208.500000 469.650000 ;
      RECT 166.500000 468.350000 199.500000 469.650000 ;
      RECT 157.500000 468.350000 158.500000 469.650000 ;
      RECT 116.500000 468.350000 149.500000 469.650000 ;
      RECT 107.500000 468.350000 108.500000 469.650000 ;
      RECT 66.500000 468.350000 99.500000 469.650000 ;
      RECT 57.500000 468.350000 58.500000 469.650000 ;
      RECT 29.500000 468.350000 49.500000 469.650000 ;
      RECT 15.500000 468.350000 16.500000 469.650000 ;
      RECT 0.000000 468.350000 2.500000 471.650000 ;
      RECT 1139.000000 467.650000 1158.500000 468.350000 ;
      RECT 732.500000 467.650000 749.000000 468.350000 ;
      RECT 666.500000 467.650000 708.500000 468.350000 ;
      RECT 616.500000 467.650000 658.500000 468.350000 ;
      RECT 566.500000 467.650000 608.500000 468.350000 ;
      RECT 516.500000 467.650000 558.500000 468.350000 ;
      RECT 466.500000 467.650000 508.500000 468.350000 ;
      RECT 416.500000 467.650000 458.500000 468.350000 ;
      RECT 366.500000 467.650000 408.500000 468.350000 ;
      RECT 316.500000 467.650000 358.500000 468.350000 ;
      RECT 266.500000 467.650000 308.500000 468.350000 ;
      RECT 216.500000 467.650000 258.500000 468.350000 ;
      RECT 166.500000 467.650000 208.500000 468.350000 ;
      RECT 116.500000 467.650000 158.500000 468.350000 ;
      RECT 66.500000 467.650000 108.500000 468.350000 ;
      RECT 29.500000 467.650000 58.500000 468.350000 ;
      RECT 0.000000 467.650000 16.500000 468.350000 ;
      RECT 1166.500000 466.350000 1186.000000 469.650000 ;
      RECT 1157.500000 466.350000 1158.500000 467.650000 ;
      RECT 732.500000 466.350000 733.500000 467.650000 ;
      RECT 716.500000 466.350000 719.500000 469.650000 ;
      RECT 707.500000 466.350000 708.500000 467.650000 ;
      RECT 666.500000 466.350000 699.500000 467.650000 ;
      RECT 657.500000 466.350000 658.500000 467.650000 ;
      RECT 616.500000 466.350000 649.500000 467.650000 ;
      RECT 607.500000 466.350000 608.500000 467.650000 ;
      RECT 566.500000 466.350000 599.500000 467.650000 ;
      RECT 557.500000 466.350000 558.500000 467.650000 ;
      RECT 516.500000 466.350000 549.500000 467.650000 ;
      RECT 507.500000 466.350000 508.500000 467.650000 ;
      RECT 466.500000 466.350000 499.500000 467.650000 ;
      RECT 457.500000 466.350000 458.500000 467.650000 ;
      RECT 416.500000 466.350000 449.500000 467.650000 ;
      RECT 407.500000 466.350000 408.500000 467.650000 ;
      RECT 366.500000 466.350000 399.500000 467.650000 ;
      RECT 357.500000 466.350000 358.500000 467.650000 ;
      RECT 316.500000 466.350000 349.500000 467.650000 ;
      RECT 307.500000 466.350000 308.500000 467.650000 ;
      RECT 266.500000 466.350000 299.500000 467.650000 ;
      RECT 257.500000 466.350000 258.500000 467.650000 ;
      RECT 216.500000 466.350000 249.500000 467.650000 ;
      RECT 207.500000 466.350000 208.500000 467.650000 ;
      RECT 166.500000 466.350000 199.500000 467.650000 ;
      RECT 157.500000 466.350000 158.500000 467.650000 ;
      RECT 116.500000 466.350000 149.500000 467.650000 ;
      RECT 107.500000 466.350000 108.500000 467.650000 ;
      RECT 66.500000 466.350000 99.500000 467.650000 ;
      RECT 57.500000 466.350000 58.500000 467.650000 ;
      RECT 29.500000 466.350000 49.500000 467.650000 ;
      RECT 15.500000 466.350000 16.500000 467.650000 ;
      RECT 1157.500000 465.650000 1186.000000 466.350000 ;
      RECT 707.500000 465.650000 733.500000 466.350000 ;
      RECT 657.500000 465.650000 699.500000 466.350000 ;
      RECT 607.500000 465.650000 649.500000 466.350000 ;
      RECT 557.500000 465.650000 599.500000 466.350000 ;
      RECT 507.500000 465.650000 549.500000 466.350000 ;
      RECT 457.500000 465.650000 499.500000 466.350000 ;
      RECT 407.500000 465.650000 449.500000 466.350000 ;
      RECT 357.500000 465.650000 399.500000 466.350000 ;
      RECT 307.500000 465.650000 349.500000 466.350000 ;
      RECT 257.500000 465.650000 299.500000 466.350000 ;
      RECT 207.500000 465.650000 249.500000 466.350000 ;
      RECT 157.500000 465.650000 199.500000 466.350000 ;
      RECT 107.500000 465.650000 149.500000 466.350000 ;
      RECT 57.500000 465.650000 99.500000 466.350000 ;
      RECT 15.500000 465.650000 49.500000 466.350000 ;
      RECT 1157.500000 464.350000 1158.500000 465.650000 ;
      RECT 1139.000000 464.350000 1149.500000 467.650000 ;
      RECT 746.500000 464.350000 749.000000 467.650000 ;
      RECT 732.500000 464.350000 733.500000 465.650000 ;
      RECT 707.500000 464.350000 708.500000 465.650000 ;
      RECT 666.500000 464.350000 699.500000 465.650000 ;
      RECT 657.500000 464.350000 658.500000 465.650000 ;
      RECT 616.500000 464.350000 649.500000 465.650000 ;
      RECT 607.500000 464.350000 608.500000 465.650000 ;
      RECT 566.500000 464.350000 599.500000 465.650000 ;
      RECT 557.500000 464.350000 558.500000 465.650000 ;
      RECT 516.500000 464.350000 549.500000 465.650000 ;
      RECT 507.500000 464.350000 508.500000 465.650000 ;
      RECT 466.500000 464.350000 499.500000 465.650000 ;
      RECT 457.500000 464.350000 458.500000 465.650000 ;
      RECT 416.500000 464.350000 449.500000 465.650000 ;
      RECT 407.500000 464.350000 408.500000 465.650000 ;
      RECT 366.500000 464.350000 399.500000 465.650000 ;
      RECT 357.500000 464.350000 358.500000 465.650000 ;
      RECT 316.500000 464.350000 349.500000 465.650000 ;
      RECT 307.500000 464.350000 308.500000 465.650000 ;
      RECT 266.500000 464.350000 299.500000 465.650000 ;
      RECT 257.500000 464.350000 258.500000 465.650000 ;
      RECT 216.500000 464.350000 249.500000 465.650000 ;
      RECT 207.500000 464.350000 208.500000 465.650000 ;
      RECT 166.500000 464.350000 199.500000 465.650000 ;
      RECT 157.500000 464.350000 158.500000 465.650000 ;
      RECT 116.500000 464.350000 149.500000 465.650000 ;
      RECT 107.500000 464.350000 108.500000 465.650000 ;
      RECT 66.500000 464.350000 99.500000 465.650000 ;
      RECT 57.500000 464.350000 58.500000 465.650000 ;
      RECT 29.500000 464.350000 49.500000 465.650000 ;
      RECT 15.500000 464.350000 16.500000 465.650000 ;
      RECT 0.000000 464.350000 2.500000 467.650000 ;
      RECT 1139.000000 463.650000 1158.500000 464.350000 ;
      RECT 732.500000 463.650000 749.000000 464.350000 ;
      RECT 666.500000 463.650000 708.500000 464.350000 ;
      RECT 616.500000 463.650000 658.500000 464.350000 ;
      RECT 566.500000 463.650000 608.500000 464.350000 ;
      RECT 516.500000 463.650000 558.500000 464.350000 ;
      RECT 466.500000 463.650000 508.500000 464.350000 ;
      RECT 416.500000 463.650000 458.500000 464.350000 ;
      RECT 366.500000 463.650000 408.500000 464.350000 ;
      RECT 316.500000 463.650000 358.500000 464.350000 ;
      RECT 266.500000 463.650000 308.500000 464.350000 ;
      RECT 216.500000 463.650000 258.500000 464.350000 ;
      RECT 166.500000 463.650000 208.500000 464.350000 ;
      RECT 116.500000 463.650000 158.500000 464.350000 ;
      RECT 66.500000 463.650000 108.500000 464.350000 ;
      RECT 29.500000 463.650000 58.500000 464.350000 ;
      RECT 0.000000 463.650000 16.500000 464.350000 ;
      RECT 1166.500000 462.350000 1186.000000 465.650000 ;
      RECT 1157.500000 462.350000 1158.500000 463.650000 ;
      RECT 732.500000 462.350000 733.500000 463.650000 ;
      RECT 716.500000 462.350000 719.500000 465.650000 ;
      RECT 707.500000 462.350000 708.500000 463.650000 ;
      RECT 666.500000 462.350000 699.500000 463.650000 ;
      RECT 657.500000 462.350000 658.500000 463.650000 ;
      RECT 616.500000 462.350000 649.500000 463.650000 ;
      RECT 607.500000 462.350000 608.500000 463.650000 ;
      RECT 566.500000 462.350000 599.500000 463.650000 ;
      RECT 557.500000 462.350000 558.500000 463.650000 ;
      RECT 516.500000 462.350000 549.500000 463.650000 ;
      RECT 507.500000 462.350000 508.500000 463.650000 ;
      RECT 466.500000 462.350000 499.500000 463.650000 ;
      RECT 457.500000 462.350000 458.500000 463.650000 ;
      RECT 416.500000 462.350000 449.500000 463.650000 ;
      RECT 407.500000 462.350000 408.500000 463.650000 ;
      RECT 366.500000 462.350000 399.500000 463.650000 ;
      RECT 357.500000 462.350000 358.500000 463.650000 ;
      RECT 316.500000 462.350000 349.500000 463.650000 ;
      RECT 307.500000 462.350000 308.500000 463.650000 ;
      RECT 266.500000 462.350000 299.500000 463.650000 ;
      RECT 257.500000 462.350000 258.500000 463.650000 ;
      RECT 216.500000 462.350000 249.500000 463.650000 ;
      RECT 207.500000 462.350000 208.500000 463.650000 ;
      RECT 166.500000 462.350000 199.500000 463.650000 ;
      RECT 157.500000 462.350000 158.500000 463.650000 ;
      RECT 116.500000 462.350000 149.500000 463.650000 ;
      RECT 107.500000 462.350000 108.500000 463.650000 ;
      RECT 66.500000 462.350000 99.500000 463.650000 ;
      RECT 57.500000 462.350000 58.500000 463.650000 ;
      RECT 29.500000 462.350000 49.500000 463.650000 ;
      RECT 15.500000 462.350000 16.500000 463.650000 ;
      RECT 1157.500000 461.650000 1186.000000 462.350000 ;
      RECT 707.500000 461.650000 733.500000 462.350000 ;
      RECT 657.500000 461.650000 699.500000 462.350000 ;
      RECT 607.500000 461.650000 649.500000 462.350000 ;
      RECT 557.500000 461.650000 599.500000 462.350000 ;
      RECT 507.500000 461.650000 549.500000 462.350000 ;
      RECT 457.500000 461.650000 499.500000 462.350000 ;
      RECT 407.500000 461.650000 449.500000 462.350000 ;
      RECT 357.500000 461.650000 399.500000 462.350000 ;
      RECT 307.500000 461.650000 349.500000 462.350000 ;
      RECT 207.500000 461.650000 249.500000 462.350000 ;
      RECT 107.500000 461.650000 149.500000 462.350000 ;
      RECT 57.500000 461.650000 99.500000 462.350000 ;
      RECT 15.500000 461.650000 49.500000 462.350000 ;
      RECT 1157.500000 460.350000 1158.500000 461.650000 ;
      RECT 1139.000000 460.350000 1149.500000 463.650000 ;
      RECT 746.500000 460.350000 749.000000 463.650000 ;
      RECT 732.500000 460.350000 733.500000 461.650000 ;
      RECT 707.500000 460.350000 708.500000 461.650000 ;
      RECT 666.500000 460.350000 699.500000 461.650000 ;
      RECT 657.500000 460.350000 658.500000 461.650000 ;
      RECT 616.500000 460.350000 649.500000 461.650000 ;
      RECT 607.500000 460.350000 608.500000 461.650000 ;
      RECT 566.500000 460.350000 599.500000 461.650000 ;
      RECT 557.500000 460.350000 558.500000 461.650000 ;
      RECT 516.500000 460.350000 549.500000 461.650000 ;
      RECT 507.500000 460.350000 508.500000 461.650000 ;
      RECT 466.500000 460.350000 499.500000 461.650000 ;
      RECT 457.500000 460.350000 458.500000 461.650000 ;
      RECT 416.500000 460.350000 449.500000 461.650000 ;
      RECT 407.500000 460.350000 408.500000 461.650000 ;
      RECT 366.500000 460.350000 399.500000 461.650000 ;
      RECT 357.500000 460.350000 358.500000 461.650000 ;
      RECT 316.500000 460.350000 349.500000 461.650000 ;
      RECT 307.500000 460.350000 308.500000 461.650000 ;
      RECT 257.500000 460.350000 299.500000 462.350000 ;
      RECT 216.500000 460.350000 249.500000 461.650000 ;
      RECT 207.500000 460.350000 208.500000 461.650000 ;
      RECT 157.500000 460.350000 199.500000 462.350000 ;
      RECT 116.500000 460.350000 149.500000 461.650000 ;
      RECT 107.500000 460.350000 108.500000 461.650000 ;
      RECT 66.500000 460.350000 99.500000 461.650000 ;
      RECT 57.500000 460.350000 58.500000 461.650000 ;
      RECT 29.500000 460.350000 49.500000 461.650000 ;
      RECT 15.500000 460.350000 16.500000 461.650000 ;
      RECT 0.000000 460.350000 2.500000 463.650000 ;
      RECT 1139.000000 459.650000 1158.500000 460.350000 ;
      RECT 732.500000 459.650000 749.000000 460.350000 ;
      RECT 666.500000 459.650000 708.500000 460.350000 ;
      RECT 616.500000 459.650000 658.500000 460.350000 ;
      RECT 566.500000 459.650000 608.500000 460.350000 ;
      RECT 516.500000 459.650000 558.500000 460.350000 ;
      RECT 466.500000 459.650000 508.500000 460.350000 ;
      RECT 416.500000 459.650000 458.500000 460.350000 ;
      RECT 366.500000 459.650000 408.500000 460.350000 ;
      RECT 316.500000 459.650000 358.500000 460.350000 ;
      RECT 216.500000 459.650000 308.500000 460.350000 ;
      RECT 116.500000 459.650000 208.500000 460.350000 ;
      RECT 66.500000 459.650000 108.500000 460.350000 ;
      RECT 29.500000 459.650000 58.500000 460.350000 ;
      RECT 0.000000 459.650000 16.500000 460.350000 ;
      RECT 1166.500000 458.350000 1186.000000 461.650000 ;
      RECT 1157.500000 458.350000 1158.500000 459.650000 ;
      RECT 732.500000 458.350000 733.500000 459.650000 ;
      RECT 716.500000 458.350000 719.500000 461.650000 ;
      RECT 707.500000 458.350000 708.500000 459.650000 ;
      RECT 666.500000 458.350000 699.500000 459.650000 ;
      RECT 657.500000 458.350000 658.500000 459.650000 ;
      RECT 616.500000 458.350000 649.500000 459.650000 ;
      RECT 607.500000 458.350000 608.500000 459.650000 ;
      RECT 566.500000 458.350000 599.500000 459.650000 ;
      RECT 557.500000 458.350000 558.500000 459.650000 ;
      RECT 516.500000 458.350000 549.500000 459.650000 ;
      RECT 507.500000 458.350000 508.500000 459.650000 ;
      RECT 466.500000 458.350000 499.500000 459.650000 ;
      RECT 457.500000 458.350000 458.500000 459.650000 ;
      RECT 416.500000 458.350000 449.500000 459.650000 ;
      RECT 407.500000 458.350000 408.500000 459.650000 ;
      RECT 366.500000 458.350000 399.500000 459.650000 ;
      RECT 357.500000 458.350000 358.500000 459.650000 ;
      RECT 316.500000 458.350000 349.500000 459.650000 ;
      RECT 307.500000 458.350000 308.500000 459.650000 ;
      RECT 216.500000 458.350000 249.500000 459.650000 ;
      RECT 207.500000 458.350000 208.500000 459.650000 ;
      RECT 116.500000 458.350000 149.500000 459.650000 ;
      RECT 107.500000 458.350000 108.500000 459.650000 ;
      RECT 66.500000 458.350000 99.500000 459.650000 ;
      RECT 57.500000 458.350000 58.500000 459.650000 ;
      RECT 29.500000 458.350000 49.500000 459.650000 ;
      RECT 15.500000 458.350000 16.500000 459.650000 ;
      RECT 1157.500000 457.650000 1186.000000 458.350000 ;
      RECT 707.500000 457.650000 733.500000 458.350000 ;
      RECT 657.500000 457.650000 699.500000 458.350000 ;
      RECT 607.500000 457.650000 649.500000 458.350000 ;
      RECT 557.500000 457.650000 599.500000 458.350000 ;
      RECT 507.500000 457.650000 549.500000 458.350000 ;
      RECT 457.500000 457.650000 499.500000 458.350000 ;
      RECT 407.500000 457.650000 449.500000 458.350000 ;
      RECT 357.500000 457.650000 399.500000 458.350000 ;
      RECT 307.500000 457.650000 349.500000 458.350000 ;
      RECT 207.500000 457.650000 249.500000 458.350000 ;
      RECT 107.500000 457.650000 149.500000 458.350000 ;
      RECT 57.500000 457.650000 99.500000 458.350000 ;
      RECT 15.500000 457.650000 49.500000 458.350000 ;
      RECT 1157.500000 456.350000 1158.500000 457.650000 ;
      RECT 1139.000000 456.350000 1149.500000 459.650000 ;
      RECT 746.500000 456.350000 749.000000 459.650000 ;
      RECT 732.500000 456.350000 733.500000 457.650000 ;
      RECT 707.500000 456.350000 708.500000 457.650000 ;
      RECT 666.500000 456.350000 699.500000 457.650000 ;
      RECT 657.500000 456.350000 658.500000 457.650000 ;
      RECT 616.500000 456.350000 649.500000 457.650000 ;
      RECT 607.500000 456.350000 608.500000 457.650000 ;
      RECT 566.500000 456.350000 599.500000 457.650000 ;
      RECT 557.500000 456.350000 558.500000 457.650000 ;
      RECT 516.500000 456.350000 549.500000 457.650000 ;
      RECT 507.500000 456.350000 508.500000 457.650000 ;
      RECT 466.500000 456.350000 499.500000 457.650000 ;
      RECT 457.500000 456.350000 458.500000 457.650000 ;
      RECT 416.500000 456.350000 449.500000 457.650000 ;
      RECT 407.500000 456.350000 408.500000 457.650000 ;
      RECT 366.500000 456.350000 399.500000 457.650000 ;
      RECT 357.500000 456.350000 358.500000 457.650000 ;
      RECT 316.500000 456.350000 349.500000 457.650000 ;
      RECT 307.500000 456.350000 308.500000 457.650000 ;
      RECT 257.500000 456.350000 299.500000 459.650000 ;
      RECT 216.500000 456.350000 249.500000 457.650000 ;
      RECT 207.500000 456.350000 208.500000 457.650000 ;
      RECT 157.500000 456.350000 199.500000 459.650000 ;
      RECT 116.500000 456.350000 149.500000 457.650000 ;
      RECT 107.500000 456.350000 108.500000 457.650000 ;
      RECT 66.500000 456.350000 99.500000 457.650000 ;
      RECT 57.500000 456.350000 58.500000 457.650000 ;
      RECT 29.500000 456.350000 49.500000 457.650000 ;
      RECT 15.500000 456.350000 16.500000 457.650000 ;
      RECT 0.000000 456.350000 2.500000 459.650000 ;
      RECT 1139.000000 455.650000 1158.500000 456.350000 ;
      RECT 732.500000 455.650000 749.000000 456.350000 ;
      RECT 666.500000 455.650000 708.500000 456.350000 ;
      RECT 616.500000 455.650000 658.500000 456.350000 ;
      RECT 566.500000 455.650000 608.500000 456.350000 ;
      RECT 516.500000 455.650000 558.500000 456.350000 ;
      RECT 466.500000 455.650000 508.500000 456.350000 ;
      RECT 416.500000 455.650000 458.500000 456.350000 ;
      RECT 366.500000 455.650000 408.500000 456.350000 ;
      RECT 316.500000 455.650000 358.500000 456.350000 ;
      RECT 216.500000 455.650000 308.500000 456.350000 ;
      RECT 116.500000 455.650000 208.500000 456.350000 ;
      RECT 66.500000 455.650000 108.500000 456.350000 ;
      RECT 29.500000 455.650000 58.500000 456.350000 ;
      RECT 0.000000 455.650000 16.500000 456.350000 ;
      RECT 1166.500000 454.350000 1186.000000 457.650000 ;
      RECT 1157.500000 454.350000 1158.500000 455.650000 ;
      RECT 732.500000 454.350000 733.500000 455.650000 ;
      RECT 716.500000 454.350000 719.500000 457.650000 ;
      RECT 707.500000 454.350000 708.500000 455.650000 ;
      RECT 666.500000 454.350000 699.500000 455.650000 ;
      RECT 657.500000 454.350000 658.500000 455.650000 ;
      RECT 616.500000 454.350000 649.500000 455.650000 ;
      RECT 607.500000 454.350000 608.500000 455.650000 ;
      RECT 566.500000 454.350000 599.500000 455.650000 ;
      RECT 557.500000 454.350000 558.500000 455.650000 ;
      RECT 516.500000 454.350000 549.500000 455.650000 ;
      RECT 507.500000 454.350000 508.500000 455.650000 ;
      RECT 466.500000 454.350000 499.500000 455.650000 ;
      RECT 457.500000 454.350000 458.500000 455.650000 ;
      RECT 416.500000 454.350000 449.500000 455.650000 ;
      RECT 407.500000 454.350000 408.500000 455.650000 ;
      RECT 366.500000 454.350000 399.500000 455.650000 ;
      RECT 357.500000 454.350000 358.500000 455.650000 ;
      RECT 316.500000 454.350000 349.500000 455.650000 ;
      RECT 307.500000 454.350000 308.500000 455.650000 ;
      RECT 216.500000 454.350000 249.500000 455.650000 ;
      RECT 207.500000 454.350000 208.500000 455.650000 ;
      RECT 116.500000 454.350000 149.500000 455.650000 ;
      RECT 107.500000 454.350000 108.500000 455.650000 ;
      RECT 66.500000 454.350000 99.500000 455.650000 ;
      RECT 57.500000 454.350000 58.500000 455.650000 ;
      RECT 29.500000 454.350000 49.500000 455.650000 ;
      RECT 15.500000 454.350000 16.500000 455.650000 ;
      RECT 1157.500000 453.650000 1186.000000 454.350000 ;
      RECT 707.500000 453.650000 733.500000 454.350000 ;
      RECT 657.500000 453.650000 699.500000 454.350000 ;
      RECT 607.500000 453.650000 649.500000 454.350000 ;
      RECT 557.500000 453.650000 599.500000 454.350000 ;
      RECT 507.500000 453.650000 549.500000 454.350000 ;
      RECT 457.500000 453.650000 499.500000 454.350000 ;
      RECT 407.500000 453.650000 449.500000 454.350000 ;
      RECT 357.500000 453.650000 399.500000 454.350000 ;
      RECT 307.500000 453.650000 349.500000 454.350000 ;
      RECT 207.500000 453.650000 249.500000 454.350000 ;
      RECT 107.500000 453.650000 149.500000 454.350000 ;
      RECT 57.500000 453.650000 99.500000 454.350000 ;
      RECT 15.500000 453.650000 49.500000 454.350000 ;
      RECT 1157.500000 452.350000 1158.500000 453.650000 ;
      RECT 1139.000000 452.350000 1149.500000 455.650000 ;
      RECT 746.500000 452.350000 749.000000 455.650000 ;
      RECT 732.500000 452.350000 733.500000 453.650000 ;
      RECT 707.500000 452.350000 708.500000 453.650000 ;
      RECT 666.500000 452.350000 699.500000 453.650000 ;
      RECT 657.500000 452.350000 658.500000 453.650000 ;
      RECT 616.500000 452.350000 649.500000 453.650000 ;
      RECT 607.500000 452.350000 608.500000 453.650000 ;
      RECT 566.500000 452.350000 599.500000 453.650000 ;
      RECT 557.500000 452.350000 558.500000 453.650000 ;
      RECT 516.500000 452.350000 549.500000 453.650000 ;
      RECT 507.500000 452.350000 508.500000 453.650000 ;
      RECT 466.500000 452.350000 499.500000 453.650000 ;
      RECT 457.500000 452.350000 458.500000 453.650000 ;
      RECT 416.500000 452.350000 449.500000 453.650000 ;
      RECT 407.500000 452.350000 408.500000 453.650000 ;
      RECT 366.500000 452.350000 399.500000 453.650000 ;
      RECT 357.500000 452.350000 358.500000 453.650000 ;
      RECT 316.500000 452.350000 349.500000 453.650000 ;
      RECT 307.500000 452.350000 308.500000 453.650000 ;
      RECT 257.500000 452.350000 299.500000 455.650000 ;
      RECT 216.500000 452.350000 249.500000 453.650000 ;
      RECT 207.500000 452.350000 208.500000 453.650000 ;
      RECT 157.500000 452.350000 199.500000 455.650000 ;
      RECT 116.500000 452.350000 149.500000 453.650000 ;
      RECT 107.500000 452.350000 108.500000 453.650000 ;
      RECT 66.500000 452.350000 99.500000 453.650000 ;
      RECT 57.500000 452.350000 58.500000 453.650000 ;
      RECT 29.500000 452.350000 49.500000 453.650000 ;
      RECT 15.500000 452.350000 16.500000 453.650000 ;
      RECT 0.000000 452.350000 2.500000 455.650000 ;
      RECT 1139.000000 451.650000 1158.500000 452.350000 ;
      RECT 732.500000 451.650000 749.000000 452.350000 ;
      RECT 666.500000 451.650000 708.500000 452.350000 ;
      RECT 616.500000 451.650000 658.500000 452.350000 ;
      RECT 566.500000 451.650000 608.500000 452.350000 ;
      RECT 516.500000 451.650000 558.500000 452.350000 ;
      RECT 466.500000 451.650000 508.500000 452.350000 ;
      RECT 416.500000 451.650000 458.500000 452.350000 ;
      RECT 366.500000 451.650000 408.500000 452.350000 ;
      RECT 316.500000 451.650000 358.500000 452.350000 ;
      RECT 216.500000 451.650000 308.500000 452.350000 ;
      RECT 116.500000 451.650000 208.500000 452.350000 ;
      RECT 66.500000 451.650000 108.500000 452.350000 ;
      RECT 29.500000 451.650000 58.500000 452.350000 ;
      RECT 0.000000 451.650000 16.500000 452.350000 ;
      RECT 1166.500000 450.350000 1186.000000 453.650000 ;
      RECT 1157.500000 450.350000 1158.500000 451.650000 ;
      RECT 732.500000 450.350000 733.500000 451.650000 ;
      RECT 716.500000 450.350000 719.500000 453.650000 ;
      RECT 707.500000 450.350000 708.500000 451.650000 ;
      RECT 666.500000 450.350000 699.500000 451.650000 ;
      RECT 657.500000 450.350000 658.500000 451.650000 ;
      RECT 616.500000 450.350000 649.500000 451.650000 ;
      RECT 607.500000 450.350000 608.500000 451.650000 ;
      RECT 566.500000 450.350000 599.500000 451.650000 ;
      RECT 557.500000 450.350000 558.500000 451.650000 ;
      RECT 516.500000 450.350000 549.500000 451.650000 ;
      RECT 507.500000 450.350000 508.500000 451.650000 ;
      RECT 466.500000 450.350000 499.500000 451.650000 ;
      RECT 457.500000 450.350000 458.500000 451.650000 ;
      RECT 416.500000 450.350000 449.500000 451.650000 ;
      RECT 407.500000 450.350000 408.500000 451.650000 ;
      RECT 366.500000 450.350000 399.500000 451.650000 ;
      RECT 357.500000 450.350000 358.500000 451.650000 ;
      RECT 316.500000 450.350000 349.500000 451.650000 ;
      RECT 307.500000 450.350000 308.500000 451.650000 ;
      RECT 216.500000 450.350000 299.500000 451.650000 ;
      RECT 207.500000 450.350000 208.500000 451.650000 ;
      RECT 116.500000 450.350000 199.500000 451.650000 ;
      RECT 107.500000 450.350000 108.500000 451.650000 ;
      RECT 66.500000 450.350000 99.500000 451.650000 ;
      RECT 57.500000 450.350000 58.500000 451.650000 ;
      RECT 29.500000 450.350000 49.500000 451.650000 ;
      RECT 15.500000 450.350000 16.500000 451.650000 ;
      RECT 1157.500000 449.650000 1186.000000 450.350000 ;
      RECT 707.500000 449.650000 733.500000 450.350000 ;
      RECT 657.500000 449.650000 699.500000 450.350000 ;
      RECT 607.500000 449.650000 649.500000 450.350000 ;
      RECT 557.500000 449.650000 599.500000 450.350000 ;
      RECT 507.500000 449.650000 549.500000 450.350000 ;
      RECT 457.500000 449.650000 499.500000 450.350000 ;
      RECT 407.500000 449.650000 449.500000 450.350000 ;
      RECT 357.500000 449.650000 399.500000 450.350000 ;
      RECT 307.500000 449.650000 349.500000 450.350000 ;
      RECT 207.500000 449.650000 299.500000 450.350000 ;
      RECT 107.500000 449.650000 199.500000 450.350000 ;
      RECT 57.500000 449.650000 99.500000 450.350000 ;
      RECT 15.500000 449.650000 49.500000 450.350000 ;
      RECT 1157.500000 448.350000 1158.500000 449.650000 ;
      RECT 1139.000000 448.350000 1149.500000 451.650000 ;
      RECT 746.500000 448.350000 749.000000 451.650000 ;
      RECT 732.500000 448.350000 733.500000 449.650000 ;
      RECT 707.500000 448.350000 708.500000 449.650000 ;
      RECT 666.500000 448.350000 699.500000 449.650000 ;
      RECT 657.500000 448.350000 658.500000 449.650000 ;
      RECT 616.500000 448.350000 649.500000 449.650000 ;
      RECT 607.500000 448.350000 608.500000 449.650000 ;
      RECT 566.500000 448.350000 599.500000 449.650000 ;
      RECT 557.500000 448.350000 558.500000 449.650000 ;
      RECT 516.500000 448.350000 549.500000 449.650000 ;
      RECT 507.500000 448.350000 508.500000 449.650000 ;
      RECT 466.500000 448.350000 499.500000 449.650000 ;
      RECT 457.500000 448.350000 458.500000 449.650000 ;
      RECT 416.500000 448.350000 449.500000 449.650000 ;
      RECT 407.500000 448.350000 408.500000 449.650000 ;
      RECT 366.500000 448.350000 399.500000 449.650000 ;
      RECT 357.500000 448.350000 358.500000 449.650000 ;
      RECT 316.500000 448.350000 349.500000 449.650000 ;
      RECT 307.500000 448.350000 308.500000 449.650000 ;
      RECT 216.500000 448.350000 299.500000 449.650000 ;
      RECT 207.500000 448.350000 208.500000 449.650000 ;
      RECT 116.500000 448.350000 199.500000 449.650000 ;
      RECT 107.500000 448.350000 108.500000 449.650000 ;
      RECT 66.500000 448.350000 99.500000 449.650000 ;
      RECT 57.500000 448.350000 58.500000 449.650000 ;
      RECT 29.500000 448.350000 49.500000 449.650000 ;
      RECT 15.500000 448.350000 16.500000 449.650000 ;
      RECT 0.000000 448.350000 2.500000 451.650000 ;
      RECT 1139.000000 447.650000 1158.500000 448.350000 ;
      RECT 732.500000 447.650000 749.000000 448.350000 ;
      RECT 666.500000 447.650000 708.500000 448.350000 ;
      RECT 616.500000 447.650000 658.500000 448.350000 ;
      RECT 566.500000 447.650000 608.500000 448.350000 ;
      RECT 516.500000 447.650000 558.500000 448.350000 ;
      RECT 466.500000 447.650000 508.500000 448.350000 ;
      RECT 416.500000 447.650000 458.500000 448.350000 ;
      RECT 366.500000 447.650000 408.500000 448.350000 ;
      RECT 316.500000 447.650000 358.500000 448.350000 ;
      RECT 216.500000 447.650000 308.500000 448.350000 ;
      RECT 116.500000 447.650000 208.500000 448.350000 ;
      RECT 66.500000 447.650000 108.500000 448.350000 ;
      RECT 29.500000 447.650000 58.500000 448.350000 ;
      RECT 0.000000 447.650000 16.500000 448.350000 ;
      RECT 1166.500000 446.350000 1186.000000 449.650000 ;
      RECT 1157.500000 446.350000 1158.500000 447.650000 ;
      RECT 732.500000 446.350000 733.500000 447.650000 ;
      RECT 716.500000 446.350000 719.500000 449.650000 ;
      RECT 707.500000 446.350000 708.500000 447.650000 ;
      RECT 666.500000 446.350000 699.500000 447.650000 ;
      RECT 657.500000 446.350000 658.500000 447.650000 ;
      RECT 616.500000 446.350000 649.500000 447.650000 ;
      RECT 607.500000 446.350000 608.500000 447.650000 ;
      RECT 566.500000 446.350000 599.500000 447.650000 ;
      RECT 557.500000 446.350000 558.500000 447.650000 ;
      RECT 516.500000 446.350000 549.500000 447.650000 ;
      RECT 507.500000 446.350000 508.500000 447.650000 ;
      RECT 466.500000 446.350000 499.500000 447.650000 ;
      RECT 457.500000 446.350000 458.500000 447.650000 ;
      RECT 416.500000 446.350000 449.500000 447.650000 ;
      RECT 407.500000 446.350000 408.500000 447.650000 ;
      RECT 366.500000 446.350000 399.500000 447.650000 ;
      RECT 357.500000 446.350000 358.500000 447.650000 ;
      RECT 316.500000 446.350000 349.500000 447.650000 ;
      RECT 307.500000 446.350000 308.500000 447.650000 ;
      RECT 216.500000 446.350000 299.500000 447.650000 ;
      RECT 207.500000 446.350000 208.500000 447.650000 ;
      RECT 116.500000 446.350000 199.500000 447.650000 ;
      RECT 107.500000 446.350000 108.500000 447.650000 ;
      RECT 66.500000 446.350000 99.500000 447.650000 ;
      RECT 57.500000 446.350000 58.500000 447.650000 ;
      RECT 29.500000 446.350000 49.500000 447.650000 ;
      RECT 15.500000 446.350000 16.500000 447.650000 ;
      RECT 1139.000000 446.000000 1149.500000 447.650000 ;
      RECT 746.500000 446.000000 749.000000 447.650000 ;
      RECT 1157.500000 445.650000 1186.000000 446.350000 ;
      RECT 746.500000 445.650000 1149.500000 446.000000 ;
      RECT 707.500000 445.650000 733.500000 446.350000 ;
      RECT 657.500000 445.650000 699.500000 446.350000 ;
      RECT 607.500000 445.650000 649.500000 446.350000 ;
      RECT 557.500000 445.650000 599.500000 446.350000 ;
      RECT 507.500000 445.650000 549.500000 446.350000 ;
      RECT 457.500000 445.650000 499.500000 446.350000 ;
      RECT 407.500000 445.650000 449.500000 446.350000 ;
      RECT 357.500000 445.650000 399.500000 446.350000 ;
      RECT 307.500000 445.650000 349.500000 446.350000 ;
      RECT 207.500000 445.650000 299.500000 446.350000 ;
      RECT 107.500000 445.650000 199.500000 446.350000 ;
      RECT 57.500000 445.650000 99.500000 446.350000 ;
      RECT 15.500000 445.650000 49.500000 446.350000 ;
      RECT 1157.500000 444.350000 1158.500000 445.650000 ;
      RECT 1116.500000 444.350000 1149.500000 445.650000 ;
      RECT 746.500000 444.350000 758.500000 445.650000 ;
      RECT 732.500000 444.350000 733.500000 445.650000 ;
      RECT 707.500000 444.350000 708.500000 445.650000 ;
      RECT 666.500000 444.350000 699.500000 445.650000 ;
      RECT 657.500000 444.350000 658.500000 445.650000 ;
      RECT 616.500000 444.350000 649.500000 445.650000 ;
      RECT 607.500000 444.350000 608.500000 445.650000 ;
      RECT 566.500000 444.350000 599.500000 445.650000 ;
      RECT 557.500000 444.350000 558.500000 445.650000 ;
      RECT 516.500000 444.350000 549.500000 445.650000 ;
      RECT 507.500000 444.350000 508.500000 445.650000 ;
      RECT 466.500000 444.350000 499.500000 445.650000 ;
      RECT 457.500000 444.350000 458.500000 445.650000 ;
      RECT 416.500000 444.350000 449.500000 445.650000 ;
      RECT 407.500000 444.350000 408.500000 445.650000 ;
      RECT 366.500000 444.350000 399.500000 445.650000 ;
      RECT 357.500000 444.350000 358.500000 445.650000 ;
      RECT 316.500000 444.350000 349.500000 445.650000 ;
      RECT 307.500000 444.350000 308.500000 445.650000 ;
      RECT 216.500000 444.350000 299.500000 445.650000 ;
      RECT 207.500000 444.350000 208.500000 445.650000 ;
      RECT 116.500000 444.350000 199.500000 445.650000 ;
      RECT 107.500000 444.350000 108.500000 445.650000 ;
      RECT 66.500000 444.350000 99.500000 445.650000 ;
      RECT 57.500000 444.350000 58.500000 445.650000 ;
      RECT 29.500000 444.350000 49.500000 445.650000 ;
      RECT 15.500000 444.350000 16.500000 445.650000 ;
      RECT 0.000000 444.350000 2.500000 447.650000 ;
      RECT 1166.500000 443.650000 1186.000000 445.650000 ;
      RECT 1116.500000 443.650000 1158.500000 444.350000 ;
      RECT 1066.500000 443.650000 1108.500000 445.650000 ;
      RECT 1016.500000 443.650000 1058.500000 445.650000 ;
      RECT 966.500000 443.650000 1008.500000 445.650000 ;
      RECT 916.500000 443.650000 958.500000 445.650000 ;
      RECT 866.500000 443.650000 908.500000 445.650000 ;
      RECT 816.500000 443.650000 858.500000 445.650000 ;
      RECT 766.500000 443.650000 808.500000 445.650000 ;
      RECT 732.500000 443.650000 758.500000 444.350000 ;
      RECT 666.500000 443.650000 708.500000 444.350000 ;
      RECT 616.500000 443.650000 658.500000 444.350000 ;
      RECT 566.500000 443.650000 608.500000 444.350000 ;
      RECT 516.500000 443.650000 558.500000 444.350000 ;
      RECT 466.500000 443.650000 508.500000 444.350000 ;
      RECT 416.500000 443.650000 458.500000 444.350000 ;
      RECT 366.500000 443.650000 408.500000 444.350000 ;
      RECT 316.500000 443.650000 358.500000 444.350000 ;
      RECT 216.500000 443.650000 308.500000 444.350000 ;
      RECT 116.500000 443.650000 208.500000 444.350000 ;
      RECT 66.500000 443.650000 108.500000 444.350000 ;
      RECT 29.500000 443.650000 58.500000 444.350000 ;
      RECT 0.000000 443.650000 16.500000 444.350000 ;
      RECT 1166.500000 442.350000 1170.500000 443.650000 ;
      RECT 1157.500000 442.350000 1158.500000 443.650000 ;
      RECT 1116.500000 442.350000 1149.500000 443.650000 ;
      RECT 1107.500000 442.350000 1108.500000 443.650000 ;
      RECT 1066.500000 442.350000 1099.500000 443.650000 ;
      RECT 1057.500000 442.350000 1058.500000 443.650000 ;
      RECT 1016.500000 442.350000 1049.500000 443.650000 ;
      RECT 1007.500000 442.350000 1008.500000 443.650000 ;
      RECT 966.500000 442.350000 999.500000 443.650000 ;
      RECT 957.500000 442.350000 958.500000 443.650000 ;
      RECT 916.500000 442.350000 949.500000 443.650000 ;
      RECT 907.500000 442.350000 908.500000 443.650000 ;
      RECT 866.500000 442.350000 899.500000 443.650000 ;
      RECT 857.500000 442.350000 858.500000 443.650000 ;
      RECT 816.500000 442.350000 849.500000 443.650000 ;
      RECT 807.500000 442.350000 808.500000 443.650000 ;
      RECT 766.500000 442.350000 799.500000 443.650000 ;
      RECT 757.500000 442.350000 758.500000 443.650000 ;
      RECT 732.500000 442.350000 733.500000 443.650000 ;
      RECT 716.500000 442.350000 719.500000 445.650000 ;
      RECT 707.500000 442.350000 708.500000 443.650000 ;
      RECT 666.500000 442.350000 699.500000 443.650000 ;
      RECT 657.500000 442.350000 658.500000 443.650000 ;
      RECT 616.500000 442.350000 649.500000 443.650000 ;
      RECT 607.500000 442.350000 608.500000 443.650000 ;
      RECT 566.500000 442.350000 599.500000 443.650000 ;
      RECT 557.500000 442.350000 558.500000 443.650000 ;
      RECT 516.500000 442.350000 549.500000 443.650000 ;
      RECT 507.500000 442.350000 508.500000 443.650000 ;
      RECT 466.500000 442.350000 499.500000 443.650000 ;
      RECT 457.500000 442.350000 458.500000 443.650000 ;
      RECT 416.500000 442.350000 449.500000 443.650000 ;
      RECT 407.500000 442.350000 408.500000 443.650000 ;
      RECT 366.500000 442.350000 399.500000 443.650000 ;
      RECT 357.500000 442.350000 358.500000 443.650000 ;
      RECT 316.500000 442.350000 349.500000 443.650000 ;
      RECT 307.500000 442.350000 308.500000 443.650000 ;
      RECT 216.500000 442.350000 299.500000 443.650000 ;
      RECT 207.500000 442.350000 208.500000 443.650000 ;
      RECT 116.500000 442.350000 199.500000 443.650000 ;
      RECT 107.500000 442.350000 108.500000 443.650000 ;
      RECT 66.500000 442.350000 99.500000 443.650000 ;
      RECT 57.500000 442.350000 58.500000 443.650000 ;
      RECT 29.500000 442.350000 49.500000 443.650000 ;
      RECT 15.500000 442.350000 16.500000 443.650000 ;
      RECT 1157.500000 441.650000 1170.500000 442.350000 ;
      RECT 1107.500000 441.650000 1149.500000 442.350000 ;
      RECT 1057.500000 441.650000 1099.500000 442.350000 ;
      RECT 1007.500000 441.650000 1049.500000 442.350000 ;
      RECT 957.500000 441.650000 999.500000 442.350000 ;
      RECT 907.500000 441.650000 949.500000 442.350000 ;
      RECT 857.500000 441.650000 899.500000 442.350000 ;
      RECT 807.500000 441.650000 849.500000 442.350000 ;
      RECT 757.500000 441.650000 799.500000 442.350000 ;
      RECT 707.500000 441.650000 733.500000 442.350000 ;
      RECT 657.500000 441.650000 699.500000 442.350000 ;
      RECT 607.500000 441.650000 649.500000 442.350000 ;
      RECT 557.500000 441.650000 599.500000 442.350000 ;
      RECT 507.500000 441.650000 549.500000 442.350000 ;
      RECT 457.500000 441.650000 499.500000 442.350000 ;
      RECT 407.500000 441.650000 449.500000 442.350000 ;
      RECT 357.500000 441.650000 399.500000 442.350000 ;
      RECT 307.500000 441.650000 349.500000 442.350000 ;
      RECT 207.500000 441.650000 299.500000 442.350000 ;
      RECT 107.500000 441.650000 199.500000 442.350000 ;
      RECT 57.500000 441.650000 99.500000 442.350000 ;
      RECT 15.500000 441.650000 49.500000 442.350000 ;
      RECT 1183.500000 440.350000 1186.000000 443.650000 ;
      RECT 1166.500000 440.350000 1170.500000 441.650000 ;
      RECT 1157.500000 440.350000 1158.500000 441.650000 ;
      RECT 1116.500000 440.350000 1149.500000 441.650000 ;
      RECT 1107.500000 440.350000 1108.500000 441.650000 ;
      RECT 1066.500000 440.350000 1099.500000 441.650000 ;
      RECT 1057.500000 440.350000 1058.500000 441.650000 ;
      RECT 1016.500000 440.350000 1049.500000 441.650000 ;
      RECT 1007.500000 440.350000 1008.500000 441.650000 ;
      RECT 966.500000 440.350000 999.500000 441.650000 ;
      RECT 957.500000 440.350000 958.500000 441.650000 ;
      RECT 916.500000 440.350000 949.500000 441.650000 ;
      RECT 907.500000 440.350000 908.500000 441.650000 ;
      RECT 866.500000 440.350000 899.500000 441.650000 ;
      RECT 857.500000 440.350000 858.500000 441.650000 ;
      RECT 816.500000 440.350000 849.500000 441.650000 ;
      RECT 807.500000 440.350000 808.500000 441.650000 ;
      RECT 766.500000 440.350000 799.500000 441.650000 ;
      RECT 757.500000 440.350000 758.500000 441.650000 ;
      RECT 746.500000 440.350000 749.500000 443.650000 ;
      RECT 732.500000 440.350000 733.500000 441.650000 ;
      RECT 707.500000 440.350000 708.500000 441.650000 ;
      RECT 666.500000 440.350000 699.500000 441.650000 ;
      RECT 657.500000 440.350000 658.500000 441.650000 ;
      RECT 616.500000 440.350000 649.500000 441.650000 ;
      RECT 607.500000 440.350000 608.500000 441.650000 ;
      RECT 566.500000 440.350000 599.500000 441.650000 ;
      RECT 557.500000 440.350000 558.500000 441.650000 ;
      RECT 516.500000 440.350000 549.500000 441.650000 ;
      RECT 507.500000 440.350000 508.500000 441.650000 ;
      RECT 466.500000 440.350000 499.500000 441.650000 ;
      RECT 457.500000 440.350000 458.500000 441.650000 ;
      RECT 416.500000 440.350000 449.500000 441.650000 ;
      RECT 407.500000 440.350000 408.500000 441.650000 ;
      RECT 366.500000 440.350000 399.500000 441.650000 ;
      RECT 357.500000 440.350000 358.500000 441.650000 ;
      RECT 316.500000 440.350000 349.500000 441.650000 ;
      RECT 307.500000 440.350000 308.500000 441.650000 ;
      RECT 216.500000 440.350000 299.500000 441.650000 ;
      RECT 207.500000 440.350000 208.500000 441.650000 ;
      RECT 116.500000 440.350000 199.500000 441.650000 ;
      RECT 107.500000 440.350000 108.500000 441.650000 ;
      RECT 66.500000 440.350000 99.500000 441.650000 ;
      RECT 57.500000 440.350000 58.500000 441.650000 ;
      RECT 29.500000 440.350000 49.500000 441.650000 ;
      RECT 15.500000 440.350000 16.500000 441.650000 ;
      RECT 0.000000 440.350000 2.500000 443.650000 ;
      RECT 1166.500000 439.650000 1186.000000 440.350000 ;
      RECT 1116.500000 439.650000 1158.500000 440.350000 ;
      RECT 1066.500000 439.650000 1108.500000 440.350000 ;
      RECT 1016.500000 439.650000 1058.500000 440.350000 ;
      RECT 966.500000 439.650000 1008.500000 440.350000 ;
      RECT 916.500000 439.650000 958.500000 440.350000 ;
      RECT 866.500000 439.650000 908.500000 440.350000 ;
      RECT 816.500000 439.650000 858.500000 440.350000 ;
      RECT 766.500000 439.650000 808.500000 440.350000 ;
      RECT 732.500000 439.650000 758.500000 440.350000 ;
      RECT 666.500000 439.650000 708.500000 440.350000 ;
      RECT 616.500000 439.650000 658.500000 440.350000 ;
      RECT 566.500000 439.650000 608.500000 440.350000 ;
      RECT 516.500000 439.650000 558.500000 440.350000 ;
      RECT 466.500000 439.650000 508.500000 440.350000 ;
      RECT 416.500000 439.650000 458.500000 440.350000 ;
      RECT 366.500000 439.650000 408.500000 440.350000 ;
      RECT 316.500000 439.650000 358.500000 440.350000 ;
      RECT 216.500000 439.650000 308.500000 440.350000 ;
      RECT 116.500000 439.650000 208.500000 440.350000 ;
      RECT 66.500000 439.650000 108.500000 440.350000 ;
      RECT 29.500000 439.650000 58.500000 440.350000 ;
      RECT 0.000000 439.650000 16.500000 440.350000 ;
      RECT 1166.500000 438.350000 1170.500000 439.650000 ;
      RECT 1157.500000 438.350000 1158.500000 439.650000 ;
      RECT 1116.500000 438.350000 1149.500000 439.650000 ;
      RECT 1107.500000 438.350000 1108.500000 439.650000 ;
      RECT 1066.500000 438.350000 1099.500000 439.650000 ;
      RECT 1057.500000 438.350000 1058.500000 439.650000 ;
      RECT 1016.500000 438.350000 1049.500000 439.650000 ;
      RECT 1007.500000 438.350000 1008.500000 439.650000 ;
      RECT 966.500000 438.350000 999.500000 439.650000 ;
      RECT 957.500000 438.350000 958.500000 439.650000 ;
      RECT 916.500000 438.350000 949.500000 439.650000 ;
      RECT 907.500000 438.350000 908.500000 439.650000 ;
      RECT 866.500000 438.350000 899.500000 439.650000 ;
      RECT 857.500000 438.350000 858.500000 439.650000 ;
      RECT 816.500000 438.350000 849.500000 439.650000 ;
      RECT 807.500000 438.350000 808.500000 439.650000 ;
      RECT 766.500000 438.350000 799.500000 439.650000 ;
      RECT 757.500000 438.350000 758.500000 439.650000 ;
      RECT 732.500000 438.350000 733.500000 439.650000 ;
      RECT 716.500000 438.350000 719.500000 441.650000 ;
      RECT 707.500000 438.350000 708.500000 439.650000 ;
      RECT 666.500000 438.350000 699.500000 439.650000 ;
      RECT 657.500000 438.350000 658.500000 439.650000 ;
      RECT 616.500000 438.350000 649.500000 439.650000 ;
      RECT 607.500000 438.350000 608.500000 439.650000 ;
      RECT 566.500000 438.350000 599.500000 439.650000 ;
      RECT 557.500000 438.350000 558.500000 439.650000 ;
      RECT 516.500000 438.350000 549.500000 439.650000 ;
      RECT 507.500000 438.350000 508.500000 439.650000 ;
      RECT 466.500000 438.350000 499.500000 439.650000 ;
      RECT 457.500000 438.350000 458.500000 439.650000 ;
      RECT 416.500000 438.350000 449.500000 439.650000 ;
      RECT 407.500000 438.350000 408.500000 439.650000 ;
      RECT 366.500000 438.350000 399.500000 439.650000 ;
      RECT 357.500000 438.350000 358.500000 439.650000 ;
      RECT 316.500000 438.350000 349.500000 439.650000 ;
      RECT 307.500000 438.350000 308.500000 439.650000 ;
      RECT 216.500000 438.350000 299.500000 439.650000 ;
      RECT 207.500000 438.350000 208.500000 439.650000 ;
      RECT 116.500000 438.350000 199.500000 439.650000 ;
      RECT 107.500000 438.350000 108.500000 439.650000 ;
      RECT 66.500000 438.350000 99.500000 439.650000 ;
      RECT 57.500000 438.350000 58.500000 439.650000 ;
      RECT 29.500000 438.350000 49.500000 439.650000 ;
      RECT 15.500000 438.350000 16.500000 439.650000 ;
      RECT 1157.500000 437.650000 1170.500000 438.350000 ;
      RECT 1107.500000 437.650000 1149.500000 438.350000 ;
      RECT 1057.500000 437.650000 1099.500000 438.350000 ;
      RECT 1007.500000 437.650000 1049.500000 438.350000 ;
      RECT 957.500000 437.650000 999.500000 438.350000 ;
      RECT 907.500000 437.650000 949.500000 438.350000 ;
      RECT 857.500000 437.650000 899.500000 438.350000 ;
      RECT 807.500000 437.650000 849.500000 438.350000 ;
      RECT 757.500000 437.650000 799.500000 438.350000 ;
      RECT 707.500000 437.650000 733.500000 438.350000 ;
      RECT 657.500000 437.650000 699.500000 438.350000 ;
      RECT 607.500000 437.650000 649.500000 438.350000 ;
      RECT 557.500000 437.650000 599.500000 438.350000 ;
      RECT 507.500000 437.650000 549.500000 438.350000 ;
      RECT 457.500000 437.650000 499.500000 438.350000 ;
      RECT 407.500000 437.650000 449.500000 438.350000 ;
      RECT 357.500000 437.650000 399.500000 438.350000 ;
      RECT 307.500000 437.650000 349.500000 438.350000 ;
      RECT 207.500000 437.650000 299.500000 438.350000 ;
      RECT 107.500000 437.650000 199.500000 438.350000 ;
      RECT 57.500000 437.650000 99.500000 438.350000 ;
      RECT 15.500000 437.650000 49.500000 438.350000 ;
      RECT 1183.500000 436.350000 1186.000000 439.650000 ;
      RECT 1166.500000 436.350000 1170.500000 437.650000 ;
      RECT 1157.500000 436.350000 1158.500000 437.650000 ;
      RECT 1116.500000 436.350000 1149.500000 437.650000 ;
      RECT 1107.500000 436.350000 1108.500000 437.650000 ;
      RECT 1066.500000 436.350000 1099.500000 437.650000 ;
      RECT 1057.500000 436.350000 1058.500000 437.650000 ;
      RECT 1016.500000 436.350000 1049.500000 437.650000 ;
      RECT 1007.500000 436.350000 1008.500000 437.650000 ;
      RECT 966.500000 436.350000 999.500000 437.650000 ;
      RECT 957.500000 436.350000 958.500000 437.650000 ;
      RECT 916.500000 436.350000 949.500000 437.650000 ;
      RECT 907.500000 436.350000 908.500000 437.650000 ;
      RECT 866.500000 436.350000 899.500000 437.650000 ;
      RECT 857.500000 436.350000 858.500000 437.650000 ;
      RECT 816.500000 436.350000 849.500000 437.650000 ;
      RECT 807.500000 436.350000 808.500000 437.650000 ;
      RECT 766.500000 436.350000 799.500000 437.650000 ;
      RECT 757.500000 436.350000 758.500000 437.650000 ;
      RECT 746.500000 436.350000 749.500000 439.650000 ;
      RECT 732.500000 436.350000 733.500000 437.650000 ;
      RECT 707.500000 436.350000 708.500000 437.650000 ;
      RECT 666.500000 436.350000 699.500000 437.650000 ;
      RECT 657.500000 436.350000 658.500000 437.650000 ;
      RECT 616.500000 436.350000 649.500000 437.650000 ;
      RECT 607.500000 436.350000 608.500000 437.650000 ;
      RECT 566.500000 436.350000 599.500000 437.650000 ;
      RECT 557.500000 436.350000 558.500000 437.650000 ;
      RECT 516.500000 436.350000 549.500000 437.650000 ;
      RECT 507.500000 436.350000 508.500000 437.650000 ;
      RECT 466.500000 436.350000 499.500000 437.650000 ;
      RECT 457.500000 436.350000 458.500000 437.650000 ;
      RECT 416.500000 436.350000 449.500000 437.650000 ;
      RECT 407.500000 436.350000 408.500000 437.650000 ;
      RECT 366.500000 436.350000 399.500000 437.650000 ;
      RECT 357.500000 436.350000 358.500000 437.650000 ;
      RECT 316.500000 436.350000 349.500000 437.650000 ;
      RECT 307.500000 436.350000 308.500000 437.650000 ;
      RECT 216.500000 436.350000 299.500000 437.650000 ;
      RECT 207.500000 436.350000 208.500000 437.650000 ;
      RECT 116.500000 436.350000 199.500000 437.650000 ;
      RECT 107.500000 436.350000 108.500000 437.650000 ;
      RECT 66.500000 436.350000 99.500000 437.650000 ;
      RECT 57.500000 436.350000 58.500000 437.650000 ;
      RECT 29.500000 436.350000 49.500000 437.650000 ;
      RECT 15.500000 436.350000 16.500000 437.650000 ;
      RECT 0.000000 436.350000 2.500000 439.650000 ;
      RECT 1166.500000 435.650000 1186.000000 436.350000 ;
      RECT 1116.500000 435.650000 1158.500000 436.350000 ;
      RECT 1066.500000 435.650000 1108.500000 436.350000 ;
      RECT 1016.500000 435.650000 1058.500000 436.350000 ;
      RECT 966.500000 435.650000 1008.500000 436.350000 ;
      RECT 916.500000 435.650000 958.500000 436.350000 ;
      RECT 866.500000 435.650000 908.500000 436.350000 ;
      RECT 816.500000 435.650000 858.500000 436.350000 ;
      RECT 766.500000 435.650000 808.500000 436.350000 ;
      RECT 732.500000 435.650000 758.500000 436.350000 ;
      RECT 666.500000 435.650000 708.500000 436.350000 ;
      RECT 616.500000 435.650000 658.500000 436.350000 ;
      RECT 566.500000 435.650000 608.500000 436.350000 ;
      RECT 516.500000 435.650000 558.500000 436.350000 ;
      RECT 466.500000 435.650000 508.500000 436.350000 ;
      RECT 416.500000 435.650000 458.500000 436.350000 ;
      RECT 366.500000 435.650000 408.500000 436.350000 ;
      RECT 316.500000 435.650000 358.500000 436.350000 ;
      RECT 216.500000 435.650000 308.500000 436.350000 ;
      RECT 116.500000 435.650000 208.500000 436.350000 ;
      RECT 66.500000 435.650000 108.500000 436.350000 ;
      RECT 29.500000 435.650000 58.500000 436.350000 ;
      RECT 0.000000 435.650000 16.500000 436.350000 ;
      RECT 1166.500000 434.350000 1170.500000 435.650000 ;
      RECT 1157.500000 434.350000 1158.500000 435.650000 ;
      RECT 1116.500000 434.350000 1149.500000 435.650000 ;
      RECT 1107.500000 434.350000 1108.500000 435.650000 ;
      RECT 1066.500000 434.350000 1099.500000 435.650000 ;
      RECT 1057.500000 434.350000 1058.500000 435.650000 ;
      RECT 1016.500000 434.350000 1049.500000 435.650000 ;
      RECT 1007.500000 434.350000 1008.500000 435.650000 ;
      RECT 966.500000 434.350000 999.500000 435.650000 ;
      RECT 957.500000 434.350000 958.500000 435.650000 ;
      RECT 916.500000 434.350000 949.500000 435.650000 ;
      RECT 907.500000 434.350000 908.500000 435.650000 ;
      RECT 866.500000 434.350000 899.500000 435.650000 ;
      RECT 857.500000 434.350000 858.500000 435.650000 ;
      RECT 816.500000 434.350000 849.500000 435.650000 ;
      RECT 807.500000 434.350000 808.500000 435.650000 ;
      RECT 766.500000 434.350000 799.500000 435.650000 ;
      RECT 757.500000 434.350000 758.500000 435.650000 ;
      RECT 732.500000 434.350000 733.500000 435.650000 ;
      RECT 716.500000 434.350000 719.500000 437.650000 ;
      RECT 707.500000 434.350000 708.500000 435.650000 ;
      RECT 666.500000 434.350000 699.500000 435.650000 ;
      RECT 657.500000 434.350000 658.500000 435.650000 ;
      RECT 616.500000 434.350000 649.500000 435.650000 ;
      RECT 607.500000 434.350000 608.500000 435.650000 ;
      RECT 566.500000 434.350000 599.500000 435.650000 ;
      RECT 557.500000 434.350000 558.500000 435.650000 ;
      RECT 516.500000 434.350000 549.500000 435.650000 ;
      RECT 507.500000 434.350000 508.500000 435.650000 ;
      RECT 466.500000 434.350000 499.500000 435.650000 ;
      RECT 457.500000 434.350000 458.500000 435.650000 ;
      RECT 416.500000 434.350000 449.500000 435.650000 ;
      RECT 407.500000 434.350000 408.500000 435.650000 ;
      RECT 366.500000 434.350000 399.500000 435.650000 ;
      RECT 357.500000 434.350000 358.500000 435.650000 ;
      RECT 316.500000 434.350000 349.500000 435.650000 ;
      RECT 307.500000 434.350000 308.500000 435.650000 ;
      RECT 216.500000 434.350000 299.500000 435.650000 ;
      RECT 207.500000 434.350000 208.500000 435.650000 ;
      RECT 116.500000 434.350000 199.500000 435.650000 ;
      RECT 107.500000 434.350000 108.500000 435.650000 ;
      RECT 66.500000 434.350000 99.500000 435.650000 ;
      RECT 57.500000 434.350000 58.500000 435.650000 ;
      RECT 29.500000 434.350000 49.500000 435.650000 ;
      RECT 15.500000 434.350000 16.500000 435.650000 ;
      RECT 1157.500000 433.650000 1170.500000 434.350000 ;
      RECT 1107.500000 433.650000 1149.500000 434.350000 ;
      RECT 1057.500000 433.650000 1099.500000 434.350000 ;
      RECT 1007.500000 433.650000 1049.500000 434.350000 ;
      RECT 957.500000 433.650000 999.500000 434.350000 ;
      RECT 907.500000 433.650000 949.500000 434.350000 ;
      RECT 857.500000 433.650000 899.500000 434.350000 ;
      RECT 807.500000 433.650000 849.500000 434.350000 ;
      RECT 757.500000 433.650000 799.500000 434.350000 ;
      RECT 707.500000 433.650000 733.500000 434.350000 ;
      RECT 657.500000 433.650000 699.500000 434.350000 ;
      RECT 607.500000 433.650000 649.500000 434.350000 ;
      RECT 557.500000 433.650000 599.500000 434.350000 ;
      RECT 507.500000 433.650000 549.500000 434.350000 ;
      RECT 457.500000 433.650000 499.500000 434.350000 ;
      RECT 407.500000 433.650000 449.500000 434.350000 ;
      RECT 357.500000 433.650000 399.500000 434.350000 ;
      RECT 307.500000 433.650000 349.500000 434.350000 ;
      RECT 207.500000 433.650000 299.500000 434.350000 ;
      RECT 107.500000 433.650000 199.500000 434.350000 ;
      RECT 57.500000 433.650000 99.500000 434.350000 ;
      RECT 15.500000 433.650000 49.500000 434.350000 ;
      RECT 1183.500000 432.350000 1186.000000 435.650000 ;
      RECT 1166.500000 432.350000 1170.500000 433.650000 ;
      RECT 1157.500000 432.350000 1158.500000 433.650000 ;
      RECT 1116.500000 432.350000 1149.500000 433.650000 ;
      RECT 1107.500000 432.350000 1108.500000 433.650000 ;
      RECT 1066.500000 432.350000 1099.500000 433.650000 ;
      RECT 1057.500000 432.350000 1058.500000 433.650000 ;
      RECT 1016.500000 432.350000 1049.500000 433.650000 ;
      RECT 1007.500000 432.350000 1008.500000 433.650000 ;
      RECT 966.500000 432.350000 999.500000 433.650000 ;
      RECT 957.500000 432.350000 958.500000 433.650000 ;
      RECT 916.500000 432.350000 949.500000 433.650000 ;
      RECT 907.500000 432.350000 908.500000 433.650000 ;
      RECT 866.500000 432.350000 899.500000 433.650000 ;
      RECT 857.500000 432.350000 858.500000 433.650000 ;
      RECT 816.500000 432.350000 849.500000 433.650000 ;
      RECT 807.500000 432.350000 808.500000 433.650000 ;
      RECT 766.500000 432.350000 799.500000 433.650000 ;
      RECT 757.500000 432.350000 758.500000 433.650000 ;
      RECT 746.500000 432.350000 749.500000 435.650000 ;
      RECT 732.500000 432.350000 733.500000 433.650000 ;
      RECT 707.500000 432.350000 708.500000 433.650000 ;
      RECT 666.500000 432.350000 699.500000 433.650000 ;
      RECT 657.500000 432.350000 658.500000 433.650000 ;
      RECT 616.500000 432.350000 649.500000 433.650000 ;
      RECT 607.500000 432.350000 608.500000 433.650000 ;
      RECT 566.500000 432.350000 599.500000 433.650000 ;
      RECT 557.500000 432.350000 558.500000 433.650000 ;
      RECT 516.500000 432.350000 549.500000 433.650000 ;
      RECT 507.500000 432.350000 508.500000 433.650000 ;
      RECT 466.500000 432.350000 499.500000 433.650000 ;
      RECT 457.500000 432.350000 458.500000 433.650000 ;
      RECT 416.500000 432.350000 449.500000 433.650000 ;
      RECT 407.500000 432.350000 408.500000 433.650000 ;
      RECT 366.500000 432.350000 399.500000 433.650000 ;
      RECT 357.500000 432.350000 358.500000 433.650000 ;
      RECT 316.500000 432.350000 349.500000 433.650000 ;
      RECT 307.500000 432.350000 308.500000 433.650000 ;
      RECT 216.500000 432.350000 299.500000 433.650000 ;
      RECT 207.500000 432.350000 208.500000 433.650000 ;
      RECT 116.500000 432.350000 199.500000 433.650000 ;
      RECT 107.500000 432.350000 108.500000 433.650000 ;
      RECT 66.500000 432.350000 99.500000 433.650000 ;
      RECT 57.500000 432.350000 58.500000 433.650000 ;
      RECT 29.500000 432.350000 49.500000 433.650000 ;
      RECT 15.500000 432.350000 16.500000 433.650000 ;
      RECT 0.000000 432.350000 2.500000 435.650000 ;
      RECT 1166.500000 431.650000 1186.000000 432.350000 ;
      RECT 1116.500000 431.650000 1158.500000 432.350000 ;
      RECT 1066.500000 431.650000 1108.500000 432.350000 ;
      RECT 1016.500000 431.650000 1058.500000 432.350000 ;
      RECT 966.500000 431.650000 1008.500000 432.350000 ;
      RECT 916.500000 431.650000 958.500000 432.350000 ;
      RECT 866.500000 431.650000 908.500000 432.350000 ;
      RECT 816.500000 431.650000 858.500000 432.350000 ;
      RECT 766.500000 431.650000 808.500000 432.350000 ;
      RECT 732.500000 431.650000 758.500000 432.350000 ;
      RECT 666.500000 431.650000 708.500000 432.350000 ;
      RECT 616.500000 431.650000 658.500000 432.350000 ;
      RECT 566.500000 431.650000 608.500000 432.350000 ;
      RECT 516.500000 431.650000 558.500000 432.350000 ;
      RECT 466.500000 431.650000 508.500000 432.350000 ;
      RECT 416.500000 431.650000 458.500000 432.350000 ;
      RECT 366.500000 431.650000 408.500000 432.350000 ;
      RECT 316.500000 431.650000 358.500000 432.350000 ;
      RECT 216.500000 431.650000 308.500000 432.350000 ;
      RECT 116.500000 431.650000 208.500000 432.350000 ;
      RECT 66.500000 431.650000 108.500000 432.350000 ;
      RECT 29.500000 431.650000 58.500000 432.350000 ;
      RECT 0.000000 431.650000 16.500000 432.350000 ;
      RECT 1166.500000 430.350000 1170.500000 431.650000 ;
      RECT 1157.500000 430.350000 1158.500000 431.650000 ;
      RECT 1116.500000 430.350000 1149.500000 431.650000 ;
      RECT 1107.500000 430.350000 1108.500000 431.650000 ;
      RECT 1066.500000 430.350000 1099.500000 431.650000 ;
      RECT 1057.500000 430.350000 1058.500000 431.650000 ;
      RECT 1016.500000 430.350000 1049.500000 431.650000 ;
      RECT 1007.500000 430.350000 1008.500000 431.650000 ;
      RECT 966.500000 430.350000 999.500000 431.650000 ;
      RECT 957.500000 430.350000 958.500000 431.650000 ;
      RECT 916.500000 430.350000 949.500000 431.650000 ;
      RECT 907.500000 430.350000 908.500000 431.650000 ;
      RECT 866.500000 430.350000 899.500000 431.650000 ;
      RECT 857.500000 430.350000 858.500000 431.650000 ;
      RECT 816.500000 430.350000 849.500000 431.650000 ;
      RECT 807.500000 430.350000 808.500000 431.650000 ;
      RECT 766.500000 430.350000 799.500000 431.650000 ;
      RECT 757.500000 430.350000 758.500000 431.650000 ;
      RECT 732.500000 430.350000 749.500000 431.650000 ;
      RECT 716.500000 430.350000 719.500000 433.650000 ;
      RECT 707.500000 430.350000 708.500000 431.650000 ;
      RECT 666.500000 430.350000 699.500000 431.650000 ;
      RECT 657.500000 430.350000 658.500000 431.650000 ;
      RECT 616.500000 430.350000 649.500000 431.650000 ;
      RECT 607.500000 430.350000 608.500000 431.650000 ;
      RECT 566.500000 430.350000 599.500000 431.650000 ;
      RECT 557.500000 430.350000 558.500000 431.650000 ;
      RECT 516.500000 430.350000 549.500000 431.650000 ;
      RECT 507.500000 430.350000 508.500000 431.650000 ;
      RECT 466.500000 430.350000 499.500000 431.650000 ;
      RECT 457.500000 430.350000 458.500000 431.650000 ;
      RECT 416.500000 430.350000 449.500000 431.650000 ;
      RECT 407.500000 430.350000 408.500000 431.650000 ;
      RECT 366.500000 430.350000 399.500000 431.650000 ;
      RECT 357.500000 430.350000 358.500000 431.650000 ;
      RECT 316.500000 430.350000 349.500000 431.650000 ;
      RECT 307.500000 430.350000 308.500000 431.650000 ;
      RECT 216.500000 430.350000 299.500000 431.650000 ;
      RECT 207.500000 430.350000 208.500000 431.650000 ;
      RECT 116.500000 430.350000 199.500000 431.650000 ;
      RECT 107.500000 430.350000 108.500000 431.650000 ;
      RECT 66.500000 430.350000 99.500000 431.650000 ;
      RECT 57.500000 430.350000 58.500000 431.650000 ;
      RECT 29.500000 430.350000 49.500000 431.650000 ;
      RECT 15.500000 430.350000 16.500000 431.650000 ;
      RECT 1157.500000 429.650000 1170.500000 430.350000 ;
      RECT 1107.500000 429.650000 1149.500000 430.350000 ;
      RECT 1057.500000 429.650000 1099.500000 430.350000 ;
      RECT 1007.500000 429.650000 1049.500000 430.350000 ;
      RECT 957.500000 429.650000 999.500000 430.350000 ;
      RECT 907.500000 429.650000 949.500000 430.350000 ;
      RECT 857.500000 429.650000 899.500000 430.350000 ;
      RECT 807.500000 429.650000 849.500000 430.350000 ;
      RECT 757.500000 429.650000 799.500000 430.350000 ;
      RECT 707.500000 429.650000 749.500000 430.350000 ;
      RECT 657.500000 429.650000 699.500000 430.350000 ;
      RECT 607.500000 429.650000 649.500000 430.350000 ;
      RECT 557.500000 429.650000 599.500000 430.350000 ;
      RECT 507.500000 429.650000 549.500000 430.350000 ;
      RECT 457.500000 429.650000 499.500000 430.350000 ;
      RECT 407.500000 429.650000 449.500000 430.350000 ;
      RECT 357.500000 429.650000 399.500000 430.350000 ;
      RECT 307.500000 429.650000 349.500000 430.350000 ;
      RECT 207.500000 429.650000 299.500000 430.350000 ;
      RECT 107.500000 429.650000 199.500000 430.350000 ;
      RECT 57.500000 429.650000 99.500000 430.350000 ;
      RECT 15.500000 429.650000 49.500000 430.350000 ;
      RECT 1183.500000 428.350000 1186.000000 431.650000 ;
      RECT 1169.500000 428.350000 1170.500000 429.650000 ;
      RECT 1116.500000 428.350000 1149.500000 429.650000 ;
      RECT 1107.500000 428.350000 1108.500000 429.650000 ;
      RECT 1066.500000 428.350000 1099.500000 429.650000 ;
      RECT 1057.500000 428.350000 1058.500000 429.650000 ;
      RECT 1016.500000 428.350000 1049.500000 429.650000 ;
      RECT 1007.500000 428.350000 1008.500000 429.650000 ;
      RECT 966.500000 428.350000 999.500000 429.650000 ;
      RECT 957.500000 428.350000 958.500000 429.650000 ;
      RECT 916.500000 428.350000 949.500000 429.650000 ;
      RECT 907.500000 428.350000 908.500000 429.650000 ;
      RECT 866.500000 428.350000 899.500000 429.650000 ;
      RECT 857.500000 428.350000 858.500000 429.650000 ;
      RECT 816.500000 428.350000 849.500000 429.650000 ;
      RECT 807.500000 428.350000 808.500000 429.650000 ;
      RECT 766.500000 428.350000 799.500000 429.650000 ;
      RECT 757.500000 428.350000 758.500000 429.650000 ;
      RECT 732.500000 428.350000 749.500000 429.650000 ;
      RECT 707.500000 428.350000 708.500000 429.650000 ;
      RECT 666.500000 428.350000 699.500000 429.650000 ;
      RECT 657.500000 428.350000 658.500000 429.650000 ;
      RECT 616.500000 428.350000 649.500000 429.650000 ;
      RECT 607.500000 428.350000 608.500000 429.650000 ;
      RECT 566.500000 428.350000 599.500000 429.650000 ;
      RECT 557.500000 428.350000 558.500000 429.650000 ;
      RECT 516.500000 428.350000 549.500000 429.650000 ;
      RECT 507.500000 428.350000 508.500000 429.650000 ;
      RECT 466.500000 428.350000 499.500000 429.650000 ;
      RECT 457.500000 428.350000 458.500000 429.650000 ;
      RECT 416.500000 428.350000 449.500000 429.650000 ;
      RECT 407.500000 428.350000 408.500000 429.650000 ;
      RECT 366.500000 428.350000 399.500000 429.650000 ;
      RECT 357.500000 428.350000 358.500000 429.650000 ;
      RECT 316.500000 428.350000 349.500000 429.650000 ;
      RECT 307.500000 428.350000 308.500000 429.650000 ;
      RECT 216.500000 428.350000 299.500000 429.650000 ;
      RECT 207.500000 428.350000 208.500000 429.650000 ;
      RECT 116.500000 428.350000 199.500000 429.650000 ;
      RECT 107.500000 428.350000 108.500000 429.650000 ;
      RECT 66.500000 428.350000 99.500000 429.650000 ;
      RECT 57.500000 428.350000 58.500000 429.650000 ;
      RECT 29.500000 428.350000 49.500000 429.650000 ;
      RECT 15.500000 428.350000 16.500000 429.650000 ;
      RECT 0.000000 428.350000 2.500000 431.650000 ;
      RECT 1169.500000 427.650000 1186.000000 428.350000 ;
      RECT 1116.500000 427.650000 1156.500000 428.350000 ;
      RECT 1066.500000 427.650000 1108.500000 428.350000 ;
      RECT 1016.500000 427.650000 1058.500000 428.350000 ;
      RECT 966.500000 427.650000 1008.500000 428.350000 ;
      RECT 916.500000 427.650000 958.500000 428.350000 ;
      RECT 866.500000 427.650000 908.500000 428.350000 ;
      RECT 816.500000 427.650000 858.500000 428.350000 ;
      RECT 766.500000 427.650000 808.500000 428.350000 ;
      RECT 732.500000 427.650000 758.500000 428.350000 ;
      RECT 666.500000 427.650000 708.500000 428.350000 ;
      RECT 616.500000 427.650000 658.500000 428.350000 ;
      RECT 566.500000 427.650000 608.500000 428.350000 ;
      RECT 516.500000 427.650000 558.500000 428.350000 ;
      RECT 466.500000 427.650000 508.500000 428.350000 ;
      RECT 416.500000 427.650000 458.500000 428.350000 ;
      RECT 366.500000 427.650000 408.500000 428.350000 ;
      RECT 316.500000 427.650000 358.500000 428.350000 ;
      RECT 216.500000 427.650000 308.500000 428.350000 ;
      RECT 116.500000 427.650000 208.500000 428.350000 ;
      RECT 66.500000 427.650000 108.500000 428.350000 ;
      RECT 29.500000 427.650000 58.500000 428.350000 ;
      RECT 0.000000 427.650000 16.500000 428.350000 ;
      RECT 1169.500000 426.350000 1170.500000 427.650000 ;
      RECT 1116.500000 426.350000 1149.500000 427.650000 ;
      RECT 1107.500000 426.350000 1108.500000 427.650000 ;
      RECT 1066.500000 426.350000 1099.500000 427.650000 ;
      RECT 1057.500000 426.350000 1058.500000 427.650000 ;
      RECT 1016.500000 426.350000 1049.500000 427.650000 ;
      RECT 1007.500000 426.350000 1008.500000 427.650000 ;
      RECT 966.500000 426.350000 999.500000 427.650000 ;
      RECT 957.500000 426.350000 958.500000 427.650000 ;
      RECT 916.500000 426.350000 949.500000 427.650000 ;
      RECT 907.500000 426.350000 908.500000 427.650000 ;
      RECT 866.500000 426.350000 899.500000 427.650000 ;
      RECT 857.500000 426.350000 858.500000 427.650000 ;
      RECT 816.500000 426.350000 849.500000 427.650000 ;
      RECT 807.500000 426.350000 808.500000 427.650000 ;
      RECT 766.500000 426.350000 799.500000 427.650000 ;
      RECT 757.500000 426.350000 758.500000 427.650000 ;
      RECT 732.500000 426.350000 749.500000 427.650000 ;
      RECT 716.500000 426.350000 719.500000 429.650000 ;
      RECT 707.500000 426.350000 708.500000 427.650000 ;
      RECT 666.500000 426.350000 699.500000 427.650000 ;
      RECT 657.500000 426.350000 658.500000 427.650000 ;
      RECT 616.500000 426.350000 649.500000 427.650000 ;
      RECT 607.500000 426.350000 608.500000 427.650000 ;
      RECT 566.500000 426.350000 599.500000 427.650000 ;
      RECT 557.500000 426.350000 558.500000 427.650000 ;
      RECT 516.500000 426.350000 549.500000 427.650000 ;
      RECT 507.500000 426.350000 508.500000 427.650000 ;
      RECT 466.500000 426.350000 499.500000 427.650000 ;
      RECT 457.500000 426.350000 458.500000 427.650000 ;
      RECT 416.500000 426.350000 449.500000 427.650000 ;
      RECT 407.500000 426.350000 408.500000 427.650000 ;
      RECT 366.500000 426.350000 399.500000 427.650000 ;
      RECT 357.500000 426.350000 358.500000 427.650000 ;
      RECT 316.500000 426.350000 349.500000 427.650000 ;
      RECT 307.500000 426.350000 308.500000 427.650000 ;
      RECT 216.500000 426.350000 299.500000 427.650000 ;
      RECT 207.500000 426.350000 208.500000 427.650000 ;
      RECT 116.500000 426.350000 199.500000 427.650000 ;
      RECT 107.500000 426.350000 108.500000 427.650000 ;
      RECT 66.500000 426.350000 99.500000 427.650000 ;
      RECT 57.500000 426.350000 58.500000 427.650000 ;
      RECT 29.500000 426.350000 49.500000 427.650000 ;
      RECT 15.500000 426.350000 16.500000 427.650000 ;
      RECT 1157.500000 425.650000 1170.500000 426.350000 ;
      RECT 1107.500000 425.650000 1149.500000 426.350000 ;
      RECT 1057.500000 425.650000 1099.500000 426.350000 ;
      RECT 1007.500000 425.650000 1049.500000 426.350000 ;
      RECT 957.500000 425.650000 999.500000 426.350000 ;
      RECT 907.500000 425.650000 949.500000 426.350000 ;
      RECT 857.500000 425.650000 899.500000 426.350000 ;
      RECT 807.500000 425.650000 849.500000 426.350000 ;
      RECT 757.500000 425.650000 799.500000 426.350000 ;
      RECT 707.500000 425.650000 749.500000 426.350000 ;
      RECT 657.500000 425.650000 699.500000 426.350000 ;
      RECT 607.500000 425.650000 649.500000 426.350000 ;
      RECT 557.500000 425.650000 599.500000 426.350000 ;
      RECT 507.500000 425.650000 549.500000 426.350000 ;
      RECT 457.500000 425.650000 499.500000 426.350000 ;
      RECT 407.500000 425.650000 449.500000 426.350000 ;
      RECT 357.500000 425.650000 399.500000 426.350000 ;
      RECT 307.500000 425.650000 349.500000 426.350000 ;
      RECT 207.500000 425.650000 299.500000 426.350000 ;
      RECT 107.500000 425.650000 199.500000 426.350000 ;
      RECT 57.500000 425.650000 99.500000 426.350000 ;
      RECT 15.500000 425.650000 49.500000 426.350000 ;
      RECT 1183.500000 424.350000 1186.000000 427.650000 ;
      RECT 1169.500000 424.350000 1170.500000 425.650000 ;
      RECT 1116.500000 424.350000 1149.500000 425.650000 ;
      RECT 1107.500000 424.350000 1108.500000 425.650000 ;
      RECT 1066.500000 424.350000 1099.500000 425.650000 ;
      RECT 1057.500000 424.350000 1058.500000 425.650000 ;
      RECT 1016.500000 424.350000 1049.500000 425.650000 ;
      RECT 1007.500000 424.350000 1008.500000 425.650000 ;
      RECT 966.500000 424.350000 999.500000 425.650000 ;
      RECT 957.500000 424.350000 958.500000 425.650000 ;
      RECT 916.500000 424.350000 949.500000 425.650000 ;
      RECT 907.500000 424.350000 908.500000 425.650000 ;
      RECT 866.500000 424.350000 899.500000 425.650000 ;
      RECT 857.500000 424.350000 858.500000 425.650000 ;
      RECT 816.500000 424.350000 849.500000 425.650000 ;
      RECT 807.500000 424.350000 808.500000 425.650000 ;
      RECT 766.500000 424.350000 799.500000 425.650000 ;
      RECT 757.500000 424.350000 758.500000 425.650000 ;
      RECT 732.500000 424.350000 749.500000 425.650000 ;
      RECT 707.500000 424.350000 708.500000 425.650000 ;
      RECT 666.500000 424.350000 699.500000 425.650000 ;
      RECT 657.500000 424.350000 658.500000 425.650000 ;
      RECT 616.500000 424.350000 649.500000 425.650000 ;
      RECT 607.500000 424.350000 608.500000 425.650000 ;
      RECT 566.500000 424.350000 599.500000 425.650000 ;
      RECT 557.500000 424.350000 558.500000 425.650000 ;
      RECT 516.500000 424.350000 549.500000 425.650000 ;
      RECT 507.500000 424.350000 508.500000 425.650000 ;
      RECT 466.500000 424.350000 499.500000 425.650000 ;
      RECT 457.500000 424.350000 458.500000 425.650000 ;
      RECT 416.500000 424.350000 449.500000 425.650000 ;
      RECT 407.500000 424.350000 408.500000 425.650000 ;
      RECT 366.500000 424.350000 399.500000 425.650000 ;
      RECT 357.500000 424.350000 358.500000 425.650000 ;
      RECT 316.500000 424.350000 349.500000 425.650000 ;
      RECT 307.500000 424.350000 308.500000 425.650000 ;
      RECT 216.500000 424.350000 299.500000 425.650000 ;
      RECT 207.500000 424.350000 208.500000 425.650000 ;
      RECT 116.500000 424.350000 199.500000 425.650000 ;
      RECT 107.500000 424.350000 108.500000 425.650000 ;
      RECT 66.500000 424.350000 99.500000 425.650000 ;
      RECT 57.500000 424.350000 58.500000 425.650000 ;
      RECT 29.500000 424.350000 49.500000 425.650000 ;
      RECT 15.500000 424.350000 16.500000 425.650000 ;
      RECT 0.000000 424.350000 2.500000 427.650000 ;
      RECT 1169.500000 423.650000 1186.000000 424.350000 ;
      RECT 1116.500000 423.650000 1156.500000 424.350000 ;
      RECT 1066.500000 423.650000 1108.500000 424.350000 ;
      RECT 1016.500000 423.650000 1058.500000 424.350000 ;
      RECT 966.500000 423.650000 1008.500000 424.350000 ;
      RECT 916.500000 423.650000 958.500000 424.350000 ;
      RECT 866.500000 423.650000 908.500000 424.350000 ;
      RECT 816.500000 423.650000 858.500000 424.350000 ;
      RECT 766.500000 423.650000 808.500000 424.350000 ;
      RECT 732.500000 423.650000 758.500000 424.350000 ;
      RECT 666.500000 423.650000 708.500000 424.350000 ;
      RECT 616.500000 423.650000 658.500000 424.350000 ;
      RECT 566.500000 423.650000 608.500000 424.350000 ;
      RECT 516.500000 423.650000 558.500000 424.350000 ;
      RECT 466.500000 423.650000 508.500000 424.350000 ;
      RECT 416.500000 423.650000 458.500000 424.350000 ;
      RECT 366.500000 423.650000 408.500000 424.350000 ;
      RECT 316.500000 423.650000 358.500000 424.350000 ;
      RECT 216.500000 423.650000 308.500000 424.350000 ;
      RECT 116.500000 423.650000 208.500000 424.350000 ;
      RECT 66.500000 423.650000 108.500000 424.350000 ;
      RECT 29.500000 423.650000 58.500000 424.350000 ;
      RECT 0.000000 423.650000 16.500000 424.350000 ;
      RECT 1169.500000 422.350000 1170.500000 423.650000 ;
      RECT 1116.500000 422.350000 1149.500000 423.650000 ;
      RECT 1107.500000 422.350000 1108.500000 423.650000 ;
      RECT 1066.500000 422.350000 1099.500000 423.650000 ;
      RECT 1057.500000 422.350000 1058.500000 423.650000 ;
      RECT 1016.500000 422.350000 1049.500000 423.650000 ;
      RECT 1007.500000 422.350000 1008.500000 423.650000 ;
      RECT 966.500000 422.350000 999.500000 423.650000 ;
      RECT 957.500000 422.350000 958.500000 423.650000 ;
      RECT 916.500000 422.350000 949.500000 423.650000 ;
      RECT 907.500000 422.350000 908.500000 423.650000 ;
      RECT 866.500000 422.350000 899.500000 423.650000 ;
      RECT 857.500000 422.350000 858.500000 423.650000 ;
      RECT 816.500000 422.350000 849.500000 423.650000 ;
      RECT 807.500000 422.350000 808.500000 423.650000 ;
      RECT 766.500000 422.350000 799.500000 423.650000 ;
      RECT 757.500000 422.350000 758.500000 423.650000 ;
      RECT 732.500000 422.350000 749.500000 423.650000 ;
      RECT 716.500000 422.350000 719.500000 425.650000 ;
      RECT 707.500000 422.350000 708.500000 423.650000 ;
      RECT 666.500000 422.350000 699.500000 423.650000 ;
      RECT 657.500000 422.350000 658.500000 423.650000 ;
      RECT 616.500000 422.350000 649.500000 423.650000 ;
      RECT 607.500000 422.350000 608.500000 423.650000 ;
      RECT 566.500000 422.350000 599.500000 423.650000 ;
      RECT 557.500000 422.350000 558.500000 423.650000 ;
      RECT 516.500000 422.350000 549.500000 423.650000 ;
      RECT 507.500000 422.350000 508.500000 423.650000 ;
      RECT 466.500000 422.350000 499.500000 423.650000 ;
      RECT 457.500000 422.350000 458.500000 423.650000 ;
      RECT 416.500000 422.350000 449.500000 423.650000 ;
      RECT 407.500000 422.350000 408.500000 423.650000 ;
      RECT 366.500000 422.350000 399.500000 423.650000 ;
      RECT 357.500000 422.350000 358.500000 423.650000 ;
      RECT 316.500000 422.350000 349.500000 423.650000 ;
      RECT 307.500000 422.350000 308.500000 423.650000 ;
      RECT 216.500000 422.350000 299.500000 423.650000 ;
      RECT 207.500000 422.350000 208.500000 423.650000 ;
      RECT 116.500000 422.350000 199.500000 423.650000 ;
      RECT 107.500000 422.350000 108.500000 423.650000 ;
      RECT 66.500000 422.350000 99.500000 423.650000 ;
      RECT 57.500000 422.350000 58.500000 423.650000 ;
      RECT 29.500000 422.350000 49.500000 423.650000 ;
      RECT 15.500000 422.350000 16.500000 423.650000 ;
      RECT 1157.500000 421.650000 1170.500000 422.350000 ;
      RECT 1107.500000 421.650000 1149.500000 422.350000 ;
      RECT 1057.500000 421.650000 1099.500000 422.350000 ;
      RECT 1007.500000 421.650000 1049.500000 422.350000 ;
      RECT 957.500000 421.650000 999.500000 422.350000 ;
      RECT 907.500000 421.650000 949.500000 422.350000 ;
      RECT 857.500000 421.650000 899.500000 422.350000 ;
      RECT 807.500000 421.650000 849.500000 422.350000 ;
      RECT 757.500000 421.650000 799.500000 422.350000 ;
      RECT 707.500000 421.650000 749.500000 422.350000 ;
      RECT 657.500000 421.650000 699.500000 422.350000 ;
      RECT 607.500000 421.650000 649.500000 422.350000 ;
      RECT 557.500000 421.650000 599.500000 422.350000 ;
      RECT 507.500000 421.650000 549.500000 422.350000 ;
      RECT 457.500000 421.650000 499.500000 422.350000 ;
      RECT 407.500000 421.650000 449.500000 422.350000 ;
      RECT 357.500000 421.650000 399.500000 422.350000 ;
      RECT 307.500000 421.650000 349.500000 422.350000 ;
      RECT 207.500000 421.650000 299.500000 422.350000 ;
      RECT 107.500000 421.650000 199.500000 422.350000 ;
      RECT 57.500000 421.650000 99.500000 422.350000 ;
      RECT 15.500000 421.650000 49.500000 422.350000 ;
      RECT 1183.500000 420.350000 1186.000000 423.650000 ;
      RECT 1169.500000 420.350000 1170.500000 421.650000 ;
      RECT 1116.500000 420.350000 1149.500000 421.650000 ;
      RECT 1107.500000 420.350000 1108.500000 421.650000 ;
      RECT 1066.500000 420.350000 1099.500000 421.650000 ;
      RECT 1057.500000 420.350000 1058.500000 421.650000 ;
      RECT 1016.500000 420.350000 1049.500000 421.650000 ;
      RECT 1007.500000 420.350000 1008.500000 421.650000 ;
      RECT 966.500000 420.350000 999.500000 421.650000 ;
      RECT 957.500000 420.350000 958.500000 421.650000 ;
      RECT 916.500000 420.350000 949.500000 421.650000 ;
      RECT 907.500000 420.350000 908.500000 421.650000 ;
      RECT 866.500000 420.350000 899.500000 421.650000 ;
      RECT 857.500000 420.350000 858.500000 421.650000 ;
      RECT 816.500000 420.350000 849.500000 421.650000 ;
      RECT 807.500000 420.350000 808.500000 421.650000 ;
      RECT 766.500000 420.350000 799.500000 421.650000 ;
      RECT 757.500000 420.350000 758.500000 421.650000 ;
      RECT 732.500000 420.350000 749.500000 421.650000 ;
      RECT 707.500000 420.350000 708.500000 421.650000 ;
      RECT 666.500000 420.350000 699.500000 421.650000 ;
      RECT 657.500000 420.350000 658.500000 421.650000 ;
      RECT 616.500000 420.350000 649.500000 421.650000 ;
      RECT 607.500000 420.350000 608.500000 421.650000 ;
      RECT 566.500000 420.350000 599.500000 421.650000 ;
      RECT 557.500000 420.350000 558.500000 421.650000 ;
      RECT 516.500000 420.350000 549.500000 421.650000 ;
      RECT 507.500000 420.350000 508.500000 421.650000 ;
      RECT 466.500000 420.350000 499.500000 421.650000 ;
      RECT 457.500000 420.350000 458.500000 421.650000 ;
      RECT 416.500000 420.350000 449.500000 421.650000 ;
      RECT 407.500000 420.350000 408.500000 421.650000 ;
      RECT 366.500000 420.350000 399.500000 421.650000 ;
      RECT 357.500000 420.350000 358.500000 421.650000 ;
      RECT 316.500000 420.350000 349.500000 421.650000 ;
      RECT 307.500000 420.350000 308.500000 421.650000 ;
      RECT 216.500000 420.350000 299.500000 421.650000 ;
      RECT 207.500000 420.350000 208.500000 421.650000 ;
      RECT 116.500000 420.350000 199.500000 421.650000 ;
      RECT 107.500000 420.350000 108.500000 421.650000 ;
      RECT 66.500000 420.350000 99.500000 421.650000 ;
      RECT 57.500000 420.350000 58.500000 421.650000 ;
      RECT 29.500000 420.350000 49.500000 421.650000 ;
      RECT 15.500000 420.350000 16.500000 421.650000 ;
      RECT 0.000000 420.350000 2.500000 423.650000 ;
      RECT 1169.500000 419.650000 1186.000000 420.350000 ;
      RECT 1116.500000 419.650000 1156.500000 420.350000 ;
      RECT 1066.500000 419.650000 1108.500000 420.350000 ;
      RECT 1016.500000 419.650000 1058.500000 420.350000 ;
      RECT 966.500000 419.650000 1008.500000 420.350000 ;
      RECT 916.500000 419.650000 958.500000 420.350000 ;
      RECT 866.500000 419.650000 908.500000 420.350000 ;
      RECT 816.500000 419.650000 858.500000 420.350000 ;
      RECT 766.500000 419.650000 808.500000 420.350000 ;
      RECT 732.500000 419.650000 758.500000 420.350000 ;
      RECT 666.500000 419.650000 708.500000 420.350000 ;
      RECT 616.500000 419.650000 658.500000 420.350000 ;
      RECT 566.500000 419.650000 608.500000 420.350000 ;
      RECT 516.500000 419.650000 558.500000 420.350000 ;
      RECT 466.500000 419.650000 508.500000 420.350000 ;
      RECT 366.500000 419.650000 408.500000 420.350000 ;
      RECT 316.500000 419.650000 358.500000 420.350000 ;
      RECT 216.500000 419.650000 308.500000 420.350000 ;
      RECT 116.500000 419.650000 208.500000 420.350000 ;
      RECT 66.500000 419.650000 108.500000 420.350000 ;
      RECT 29.500000 419.650000 58.500000 420.350000 ;
      RECT 0.000000 419.650000 16.500000 420.350000 ;
      RECT 416.500000 418.605000 458.500000 420.350000 ;
      RECT 1169.500000 418.350000 1170.500000 419.650000 ;
      RECT 1116.500000 418.350000 1149.500000 419.650000 ;
      RECT 1107.500000 418.350000 1108.500000 419.650000 ;
      RECT 1066.500000 418.350000 1099.500000 419.650000 ;
      RECT 1057.500000 418.350000 1058.500000 419.650000 ;
      RECT 1016.500000 418.350000 1049.500000 419.650000 ;
      RECT 1007.500000 418.350000 1008.500000 419.650000 ;
      RECT 966.500000 418.350000 999.500000 419.650000 ;
      RECT 957.500000 418.350000 958.500000 419.650000 ;
      RECT 916.500000 418.350000 949.500000 419.650000 ;
      RECT 907.500000 418.350000 908.500000 419.650000 ;
      RECT 866.500000 418.350000 899.500000 419.650000 ;
      RECT 857.500000 418.350000 858.500000 419.650000 ;
      RECT 816.500000 418.350000 849.500000 419.650000 ;
      RECT 807.500000 418.350000 808.500000 419.650000 ;
      RECT 766.500000 418.350000 799.500000 419.650000 ;
      RECT 757.500000 418.350000 758.500000 419.650000 ;
      RECT 732.500000 418.350000 749.500000 419.650000 ;
      RECT 716.500000 418.350000 719.500000 421.650000 ;
      RECT 707.500000 418.350000 708.500000 419.650000 ;
      RECT 666.500000 418.350000 699.500000 419.650000 ;
      RECT 657.500000 418.350000 658.500000 419.650000 ;
      RECT 616.500000 418.350000 649.500000 419.650000 ;
      RECT 607.500000 418.350000 608.500000 419.650000 ;
      RECT 566.500000 418.350000 599.500000 419.650000 ;
      RECT 557.500000 418.350000 558.500000 419.650000 ;
      RECT 516.500000 418.350000 549.500000 419.650000 ;
      RECT 507.500000 418.350000 508.500000 419.650000 ;
      RECT 466.500000 418.350000 499.500000 419.650000 ;
      RECT 457.500000 418.350000 458.500000 418.605000 ;
      RECT 416.500000 418.350000 449.500000 418.605000 ;
      RECT 407.500000 418.350000 408.500000 419.650000 ;
      RECT 366.500000 418.350000 399.500000 419.650000 ;
      RECT 357.500000 418.350000 358.500000 419.650000 ;
      RECT 316.500000 418.350000 349.500000 419.650000 ;
      RECT 307.500000 418.350000 308.500000 419.650000 ;
      RECT 216.500000 418.350000 299.500000 419.650000 ;
      RECT 207.500000 418.350000 208.500000 419.650000 ;
      RECT 116.500000 418.350000 199.500000 419.650000 ;
      RECT 107.500000 418.350000 108.500000 419.650000 ;
      RECT 66.500000 418.350000 99.500000 419.650000 ;
      RECT 57.500000 418.350000 58.500000 419.650000 ;
      RECT 29.500000 418.350000 49.500000 419.650000 ;
      RECT 15.500000 418.350000 16.500000 419.650000 ;
      RECT 1157.500000 417.650000 1170.500000 418.350000 ;
      RECT 1107.500000 417.650000 1149.500000 418.350000 ;
      RECT 1057.500000 417.650000 1099.500000 418.350000 ;
      RECT 1007.500000 417.650000 1049.500000 418.350000 ;
      RECT 957.500000 417.650000 999.500000 418.350000 ;
      RECT 907.500000 417.650000 949.500000 418.350000 ;
      RECT 857.500000 417.650000 899.500000 418.350000 ;
      RECT 807.500000 417.650000 849.500000 418.350000 ;
      RECT 757.500000 417.650000 799.500000 418.350000 ;
      RECT 707.500000 417.650000 749.500000 418.350000 ;
      RECT 657.500000 417.650000 699.500000 418.350000 ;
      RECT 607.500000 417.650000 649.500000 418.350000 ;
      RECT 557.500000 417.650000 599.500000 418.350000 ;
      RECT 507.500000 417.650000 549.500000 418.350000 ;
      RECT 407.500000 417.650000 449.500000 418.350000 ;
      RECT 357.500000 417.650000 399.500000 418.350000 ;
      RECT 307.500000 417.650000 349.500000 418.350000 ;
      RECT 207.500000 417.650000 299.500000 418.350000 ;
      RECT 107.500000 417.650000 199.500000 418.350000 ;
      RECT 57.500000 417.650000 99.500000 418.350000 ;
      RECT 15.500000 417.650000 49.500000 418.350000 ;
      RECT 1183.500000 416.350000 1186.000000 419.650000 ;
      RECT 1169.500000 416.350000 1170.500000 417.650000 ;
      RECT 1116.500000 416.350000 1149.500000 417.650000 ;
      RECT 1107.500000 416.350000 1108.500000 417.650000 ;
      RECT 1066.500000 416.350000 1099.500000 417.650000 ;
      RECT 1057.500000 416.350000 1058.500000 417.650000 ;
      RECT 1016.500000 416.350000 1049.500000 417.650000 ;
      RECT 1007.500000 416.350000 1008.500000 417.650000 ;
      RECT 966.500000 416.350000 999.500000 417.650000 ;
      RECT 957.500000 416.350000 958.500000 417.650000 ;
      RECT 916.500000 416.350000 949.500000 417.650000 ;
      RECT 907.500000 416.350000 908.500000 417.650000 ;
      RECT 866.500000 416.350000 899.500000 417.650000 ;
      RECT 857.500000 416.350000 858.500000 417.650000 ;
      RECT 816.500000 416.350000 849.500000 417.650000 ;
      RECT 807.500000 416.350000 808.500000 417.650000 ;
      RECT 766.500000 416.350000 799.500000 417.650000 ;
      RECT 757.500000 416.350000 758.500000 417.650000 ;
      RECT 716.500000 416.350000 749.500000 417.650000 ;
      RECT 707.500000 416.350000 708.500000 417.650000 ;
      RECT 666.500000 416.350000 699.500000 417.650000 ;
      RECT 657.500000 416.350000 658.500000 417.650000 ;
      RECT 616.500000 416.350000 649.500000 417.650000 ;
      RECT 607.500000 416.350000 608.500000 417.650000 ;
      RECT 566.500000 416.350000 599.500000 417.650000 ;
      RECT 557.500000 416.350000 558.500000 417.650000 ;
      RECT 516.500000 416.350000 549.500000 417.650000 ;
      RECT 507.500000 416.350000 508.500000 417.650000 ;
      RECT 457.500000 416.350000 499.500000 418.350000 ;
      RECT 407.500000 416.350000 408.500000 417.650000 ;
      RECT 366.500000 416.350000 399.500000 417.650000 ;
      RECT 357.500000 416.350000 358.500000 417.650000 ;
      RECT 316.500000 416.350000 349.500000 417.650000 ;
      RECT 307.500000 416.350000 308.500000 417.650000 ;
      RECT 216.500000 416.350000 299.500000 417.650000 ;
      RECT 207.500000 416.350000 208.500000 417.650000 ;
      RECT 116.500000 416.350000 199.500000 417.650000 ;
      RECT 107.500000 416.350000 108.500000 417.650000 ;
      RECT 66.500000 416.350000 99.500000 417.650000 ;
      RECT 57.500000 416.350000 58.500000 417.650000 ;
      RECT 29.500000 416.350000 49.500000 417.650000 ;
      RECT 15.500000 416.350000 16.500000 417.650000 ;
      RECT 0.000000 416.350000 2.500000 419.650000 ;
      RECT 1169.500000 415.650000 1186.000000 416.350000 ;
      RECT 1116.500000 415.650000 1156.500000 416.350000 ;
      RECT 1066.500000 415.650000 1108.500000 416.350000 ;
      RECT 1016.500000 415.650000 1058.500000 416.350000 ;
      RECT 966.500000 415.650000 1008.500000 416.350000 ;
      RECT 916.500000 415.650000 958.500000 416.350000 ;
      RECT 866.500000 415.650000 908.500000 416.350000 ;
      RECT 816.500000 415.650000 858.500000 416.350000 ;
      RECT 766.500000 415.650000 808.500000 416.350000 ;
      RECT 716.500000 415.650000 758.500000 416.350000 ;
      RECT 666.500000 415.650000 708.500000 416.350000 ;
      RECT 616.500000 415.650000 658.500000 416.350000 ;
      RECT 566.500000 415.650000 608.500000 416.350000 ;
      RECT 516.500000 415.650000 558.500000 416.350000 ;
      RECT 457.500000 415.650000 508.500000 416.350000 ;
      RECT 366.500000 415.650000 408.500000 416.350000 ;
      RECT 316.500000 415.650000 358.500000 416.350000 ;
      RECT 216.500000 415.650000 308.500000 416.350000 ;
      RECT 116.500000 415.650000 208.500000 416.350000 ;
      RECT 66.500000 415.650000 108.500000 416.350000 ;
      RECT 29.500000 415.650000 58.500000 416.350000 ;
      RECT 0.000000 415.650000 16.500000 416.350000 ;
      RECT 457.500000 414.605000 499.500000 415.650000 ;
      RECT 416.500000 414.605000 449.500000 417.650000 ;
      RECT 1169.500000 414.350000 1170.500000 415.650000 ;
      RECT 1116.500000 414.350000 1149.500000 415.650000 ;
      RECT 1107.500000 414.350000 1108.500000 415.650000 ;
      RECT 1066.500000 414.350000 1099.500000 415.650000 ;
      RECT 1057.500000 414.350000 1058.500000 415.650000 ;
      RECT 1016.500000 414.350000 1049.500000 415.650000 ;
      RECT 1007.500000 414.350000 1008.500000 415.650000 ;
      RECT 966.500000 414.350000 999.500000 415.650000 ;
      RECT 957.500000 414.350000 958.500000 415.650000 ;
      RECT 916.500000 414.350000 949.500000 415.650000 ;
      RECT 907.500000 414.350000 908.500000 415.650000 ;
      RECT 866.500000 414.350000 899.500000 415.650000 ;
      RECT 857.500000 414.350000 858.500000 415.650000 ;
      RECT 816.500000 414.350000 849.500000 415.650000 ;
      RECT 807.500000 414.350000 808.500000 415.650000 ;
      RECT 766.500000 414.350000 799.500000 415.650000 ;
      RECT 757.500000 414.350000 758.500000 415.650000 ;
      RECT 716.500000 414.350000 749.500000 415.650000 ;
      RECT 707.500000 414.350000 708.500000 415.650000 ;
      RECT 666.500000 414.350000 699.500000 415.650000 ;
      RECT 657.500000 414.350000 658.500000 415.650000 ;
      RECT 616.500000 414.350000 649.500000 415.650000 ;
      RECT 607.500000 414.350000 608.500000 415.650000 ;
      RECT 566.500000 414.350000 599.500000 415.650000 ;
      RECT 557.500000 414.350000 558.500000 415.650000 ;
      RECT 516.500000 414.350000 549.500000 415.650000 ;
      RECT 507.500000 414.350000 508.500000 415.650000 ;
      RECT 416.500000 414.350000 499.500000 414.605000 ;
      RECT 407.500000 414.350000 408.500000 415.650000 ;
      RECT 366.500000 414.350000 399.500000 415.650000 ;
      RECT 357.500000 414.350000 358.500000 415.650000 ;
      RECT 316.500000 414.350000 349.500000 415.650000 ;
      RECT 307.500000 414.350000 308.500000 415.650000 ;
      RECT 216.500000 414.350000 299.500000 415.650000 ;
      RECT 207.500000 414.350000 208.500000 415.650000 ;
      RECT 116.500000 414.350000 199.500000 415.650000 ;
      RECT 107.500000 414.350000 108.500000 415.650000 ;
      RECT 66.500000 414.350000 99.500000 415.650000 ;
      RECT 57.500000 414.350000 58.500000 415.650000 ;
      RECT 29.500000 414.350000 49.500000 415.650000 ;
      RECT 15.500000 414.350000 16.500000 415.650000 ;
      RECT 1157.500000 413.650000 1170.500000 414.350000 ;
      RECT 1107.500000 413.650000 1149.500000 414.350000 ;
      RECT 1057.500000 413.650000 1099.500000 414.350000 ;
      RECT 1007.500000 413.650000 1049.500000 414.350000 ;
      RECT 957.500000 413.650000 999.500000 414.350000 ;
      RECT 907.500000 413.650000 949.500000 414.350000 ;
      RECT 857.500000 413.650000 899.500000 414.350000 ;
      RECT 807.500000 413.650000 849.500000 414.350000 ;
      RECT 757.500000 413.650000 799.500000 414.350000 ;
      RECT 707.500000 413.650000 749.500000 414.350000 ;
      RECT 657.500000 413.650000 699.500000 414.350000 ;
      RECT 607.500000 413.650000 649.500000 414.350000 ;
      RECT 557.500000 413.650000 599.500000 414.350000 ;
      RECT 507.500000 413.650000 549.500000 414.350000 ;
      RECT 407.500000 413.650000 499.500000 414.350000 ;
      RECT 357.500000 413.650000 399.500000 414.350000 ;
      RECT 307.500000 413.650000 349.500000 414.350000 ;
      RECT 207.500000 413.650000 299.500000 414.350000 ;
      RECT 107.500000 413.650000 199.500000 414.350000 ;
      RECT 57.500000 413.650000 99.500000 414.350000 ;
      RECT 15.500000 413.650000 49.500000 414.350000 ;
      RECT 1183.500000 412.350000 1186.000000 415.650000 ;
      RECT 1169.500000 412.350000 1170.500000 413.650000 ;
      RECT 1116.500000 412.350000 1149.500000 413.650000 ;
      RECT 1107.500000 412.350000 1108.500000 413.650000 ;
      RECT 1066.500000 412.350000 1099.500000 413.650000 ;
      RECT 1057.500000 412.350000 1058.500000 413.650000 ;
      RECT 1016.500000 412.350000 1049.500000 413.650000 ;
      RECT 1007.500000 412.350000 1008.500000 413.650000 ;
      RECT 966.500000 412.350000 999.500000 413.650000 ;
      RECT 957.500000 412.350000 958.500000 413.650000 ;
      RECT 916.500000 412.350000 949.500000 413.650000 ;
      RECT 907.500000 412.350000 908.500000 413.650000 ;
      RECT 866.500000 412.350000 899.500000 413.650000 ;
      RECT 857.500000 412.350000 858.500000 413.650000 ;
      RECT 816.500000 412.350000 849.500000 413.650000 ;
      RECT 807.500000 412.350000 808.500000 413.650000 ;
      RECT 766.500000 412.350000 799.500000 413.650000 ;
      RECT 757.500000 412.350000 758.500000 413.650000 ;
      RECT 716.500000 412.350000 749.500000 413.650000 ;
      RECT 707.500000 412.350000 708.500000 413.650000 ;
      RECT 666.500000 412.350000 699.500000 413.650000 ;
      RECT 657.500000 412.350000 658.500000 413.650000 ;
      RECT 616.500000 412.350000 649.500000 413.650000 ;
      RECT 607.500000 412.350000 608.500000 413.650000 ;
      RECT 566.500000 412.350000 599.500000 413.650000 ;
      RECT 557.500000 412.350000 558.500000 413.650000 ;
      RECT 516.500000 412.350000 549.500000 413.650000 ;
      RECT 507.500000 412.350000 508.500000 413.650000 ;
      RECT 416.500000 412.350000 499.500000 413.650000 ;
      RECT 407.500000 412.350000 408.500000 413.650000 ;
      RECT 366.500000 412.350000 399.500000 413.650000 ;
      RECT 357.500000 412.350000 358.500000 413.650000 ;
      RECT 316.500000 412.350000 349.500000 413.650000 ;
      RECT 307.500000 412.350000 308.500000 413.650000 ;
      RECT 216.500000 412.350000 299.500000 413.650000 ;
      RECT 207.500000 412.350000 208.500000 413.650000 ;
      RECT 116.500000 412.350000 199.500000 413.650000 ;
      RECT 107.500000 412.350000 108.500000 413.650000 ;
      RECT 66.500000 412.350000 99.500000 413.650000 ;
      RECT 57.500000 412.350000 58.500000 413.650000 ;
      RECT 29.500000 412.350000 49.500000 413.650000 ;
      RECT 15.500000 412.350000 16.500000 413.650000 ;
      RECT 0.000000 412.350000 2.500000 415.650000 ;
      RECT 1169.500000 411.650000 1186.000000 412.350000 ;
      RECT 1116.500000 411.650000 1156.500000 412.350000 ;
      RECT 1066.500000 411.650000 1108.500000 412.350000 ;
      RECT 1016.500000 411.650000 1058.500000 412.350000 ;
      RECT 966.500000 411.650000 1008.500000 412.350000 ;
      RECT 916.500000 411.650000 958.500000 412.350000 ;
      RECT 866.500000 411.650000 908.500000 412.350000 ;
      RECT 816.500000 411.650000 858.500000 412.350000 ;
      RECT 766.500000 411.650000 808.500000 412.350000 ;
      RECT 716.500000 411.650000 758.500000 412.350000 ;
      RECT 666.500000 411.650000 708.500000 412.350000 ;
      RECT 616.500000 411.650000 658.500000 412.350000 ;
      RECT 566.500000 411.650000 608.500000 412.350000 ;
      RECT 516.500000 411.650000 558.500000 412.350000 ;
      RECT 416.500000 411.650000 508.500000 412.350000 ;
      RECT 366.500000 411.650000 408.500000 412.350000 ;
      RECT 316.500000 411.650000 358.500000 412.350000 ;
      RECT 216.500000 411.650000 308.500000 412.350000 ;
      RECT 116.500000 411.650000 208.500000 412.350000 ;
      RECT 66.500000 411.650000 108.500000 412.350000 ;
      RECT 29.500000 411.650000 58.500000 412.350000 ;
      RECT 0.000000 411.650000 16.500000 412.350000 ;
      RECT 1169.500000 410.350000 1170.500000 411.650000 ;
      RECT 1116.500000 410.350000 1149.500000 411.650000 ;
      RECT 1107.500000 410.350000 1108.500000 411.650000 ;
      RECT 1066.500000 410.350000 1099.500000 411.650000 ;
      RECT 1057.500000 410.350000 1058.500000 411.650000 ;
      RECT 1016.500000 410.350000 1049.500000 411.650000 ;
      RECT 1007.500000 410.350000 1008.500000 411.650000 ;
      RECT 966.500000 410.350000 999.500000 411.650000 ;
      RECT 957.500000 410.350000 958.500000 411.650000 ;
      RECT 916.500000 410.350000 949.500000 411.650000 ;
      RECT 907.500000 410.350000 908.500000 411.650000 ;
      RECT 866.500000 410.350000 899.500000 411.650000 ;
      RECT 857.500000 410.350000 858.500000 411.650000 ;
      RECT 816.500000 410.350000 849.500000 411.650000 ;
      RECT 807.500000 410.350000 808.500000 411.650000 ;
      RECT 766.500000 410.350000 799.500000 411.650000 ;
      RECT 757.500000 410.350000 758.500000 411.650000 ;
      RECT 716.500000 410.350000 749.500000 411.650000 ;
      RECT 707.500000 410.350000 708.500000 411.650000 ;
      RECT 666.500000 410.350000 699.500000 411.650000 ;
      RECT 657.500000 410.350000 658.500000 411.650000 ;
      RECT 616.500000 410.350000 649.500000 411.650000 ;
      RECT 607.500000 410.350000 608.500000 411.650000 ;
      RECT 566.500000 410.350000 599.500000 411.650000 ;
      RECT 557.500000 410.350000 558.500000 411.650000 ;
      RECT 516.500000 410.350000 549.500000 411.650000 ;
      RECT 507.500000 410.350000 508.500000 411.650000 ;
      RECT 416.500000 410.350000 499.500000 411.650000 ;
      RECT 407.500000 410.350000 408.500000 411.650000 ;
      RECT 366.500000 410.350000 399.500000 411.650000 ;
      RECT 357.500000 410.350000 358.500000 411.650000 ;
      RECT 316.500000 410.350000 349.500000 411.650000 ;
      RECT 307.500000 410.350000 308.500000 411.650000 ;
      RECT 216.500000 410.350000 299.500000 411.650000 ;
      RECT 207.500000 410.350000 208.500000 411.650000 ;
      RECT 116.500000 410.350000 199.500000 411.650000 ;
      RECT 107.500000 410.350000 108.500000 411.650000 ;
      RECT 66.500000 410.350000 99.500000 411.650000 ;
      RECT 57.500000 410.350000 58.500000 411.650000 ;
      RECT 29.500000 410.350000 49.500000 411.650000 ;
      RECT 15.500000 410.350000 16.500000 411.650000 ;
      RECT 1157.500000 409.650000 1170.500000 410.350000 ;
      RECT 1107.500000 409.650000 1149.500000 410.350000 ;
      RECT 1057.500000 409.650000 1099.500000 410.350000 ;
      RECT 1007.500000 409.650000 1049.500000 410.350000 ;
      RECT 957.500000 409.650000 999.500000 410.350000 ;
      RECT 907.500000 409.650000 949.500000 410.350000 ;
      RECT 857.500000 409.650000 899.500000 410.350000 ;
      RECT 807.500000 409.650000 849.500000 410.350000 ;
      RECT 757.500000 409.650000 799.500000 410.350000 ;
      RECT 707.500000 409.650000 749.500000 410.350000 ;
      RECT 657.500000 409.650000 699.500000 410.350000 ;
      RECT 607.500000 409.650000 649.500000 410.350000 ;
      RECT 557.500000 409.650000 599.500000 410.350000 ;
      RECT 507.500000 409.650000 549.500000 410.350000 ;
      RECT 407.500000 409.650000 499.500000 410.350000 ;
      RECT 357.500000 409.650000 399.500000 410.350000 ;
      RECT 307.500000 409.650000 349.500000 410.350000 ;
      RECT 207.500000 409.650000 299.500000 410.350000 ;
      RECT 107.500000 409.650000 199.500000 410.350000 ;
      RECT 57.500000 409.650000 99.500000 410.350000 ;
      RECT 15.500000 409.650000 49.500000 410.350000 ;
      RECT 1183.500000 408.350000 1186.000000 411.650000 ;
      RECT 1169.500000 408.350000 1170.500000 409.650000 ;
      RECT 1116.500000 408.350000 1149.500000 409.650000 ;
      RECT 1107.500000 408.350000 1108.500000 409.650000 ;
      RECT 1066.500000 408.350000 1099.500000 409.650000 ;
      RECT 1057.500000 408.350000 1058.500000 409.650000 ;
      RECT 1016.500000 408.350000 1049.500000 409.650000 ;
      RECT 1007.500000 408.350000 1008.500000 409.650000 ;
      RECT 966.500000 408.350000 999.500000 409.650000 ;
      RECT 957.500000 408.350000 958.500000 409.650000 ;
      RECT 916.500000 408.350000 949.500000 409.650000 ;
      RECT 907.500000 408.350000 908.500000 409.650000 ;
      RECT 866.500000 408.350000 899.500000 409.650000 ;
      RECT 857.500000 408.350000 858.500000 409.650000 ;
      RECT 816.500000 408.350000 849.500000 409.650000 ;
      RECT 807.500000 408.350000 808.500000 409.650000 ;
      RECT 766.500000 408.350000 799.500000 409.650000 ;
      RECT 757.500000 408.350000 758.500000 409.650000 ;
      RECT 716.500000 408.350000 749.500000 409.650000 ;
      RECT 707.500000 408.350000 708.500000 409.650000 ;
      RECT 666.500000 408.350000 699.500000 409.650000 ;
      RECT 657.500000 408.350000 658.500000 409.650000 ;
      RECT 616.500000 408.350000 649.500000 409.650000 ;
      RECT 607.500000 408.350000 608.500000 409.650000 ;
      RECT 566.500000 408.350000 599.500000 409.650000 ;
      RECT 557.500000 408.350000 558.500000 409.650000 ;
      RECT 516.500000 408.350000 549.500000 409.650000 ;
      RECT 507.500000 408.350000 508.500000 409.650000 ;
      RECT 416.500000 408.350000 499.500000 409.650000 ;
      RECT 407.500000 408.350000 408.500000 409.650000 ;
      RECT 366.500000 408.350000 399.500000 409.650000 ;
      RECT 357.500000 408.350000 358.500000 409.650000 ;
      RECT 316.500000 408.350000 349.500000 409.650000 ;
      RECT 307.500000 408.350000 308.500000 409.650000 ;
      RECT 216.500000 408.350000 299.500000 409.650000 ;
      RECT 207.500000 408.350000 208.500000 409.650000 ;
      RECT 116.500000 408.350000 199.500000 409.650000 ;
      RECT 107.500000 408.350000 108.500000 409.650000 ;
      RECT 66.500000 408.350000 99.500000 409.650000 ;
      RECT 57.500000 408.350000 58.500000 409.650000 ;
      RECT 29.500000 408.350000 49.500000 409.650000 ;
      RECT 15.500000 408.350000 16.500000 409.650000 ;
      RECT 0.000000 408.350000 2.500000 411.650000 ;
      RECT 1169.500000 407.650000 1186.000000 408.350000 ;
      RECT 1116.500000 407.650000 1156.500000 408.350000 ;
      RECT 1066.500000 407.650000 1108.500000 408.350000 ;
      RECT 1016.500000 407.650000 1058.500000 408.350000 ;
      RECT 966.500000 407.650000 1008.500000 408.350000 ;
      RECT 916.500000 407.650000 958.500000 408.350000 ;
      RECT 866.500000 407.650000 908.500000 408.350000 ;
      RECT 816.500000 407.650000 858.500000 408.350000 ;
      RECT 766.500000 407.650000 808.500000 408.350000 ;
      RECT 716.500000 407.650000 758.500000 408.350000 ;
      RECT 666.500000 407.650000 708.500000 408.350000 ;
      RECT 616.500000 407.650000 658.500000 408.350000 ;
      RECT 566.500000 407.650000 608.500000 408.350000 ;
      RECT 516.500000 407.650000 558.500000 408.350000 ;
      RECT 416.500000 407.650000 508.500000 408.350000 ;
      RECT 366.500000 407.650000 408.500000 408.350000 ;
      RECT 316.500000 407.650000 358.500000 408.350000 ;
      RECT 216.500000 407.650000 308.500000 408.350000 ;
      RECT 116.500000 407.650000 208.500000 408.350000 ;
      RECT 66.500000 407.650000 108.500000 408.350000 ;
      RECT 29.500000 407.650000 58.500000 408.350000 ;
      RECT 0.000000 407.650000 16.500000 408.350000 ;
      RECT 1169.500000 406.350000 1170.500000 407.650000 ;
      RECT 1116.500000 406.350000 1149.500000 407.650000 ;
      RECT 1107.500000 406.350000 1108.500000 407.650000 ;
      RECT 1066.500000 406.350000 1099.500000 407.650000 ;
      RECT 1057.500000 406.350000 1058.500000 407.650000 ;
      RECT 1016.500000 406.350000 1049.500000 407.650000 ;
      RECT 1007.500000 406.350000 1008.500000 407.650000 ;
      RECT 966.500000 406.350000 999.500000 407.650000 ;
      RECT 957.500000 406.350000 958.500000 407.650000 ;
      RECT 916.500000 406.350000 949.500000 407.650000 ;
      RECT 907.500000 406.350000 908.500000 407.650000 ;
      RECT 866.500000 406.350000 899.500000 407.650000 ;
      RECT 857.500000 406.350000 858.500000 407.650000 ;
      RECT 816.500000 406.350000 849.500000 407.650000 ;
      RECT 807.500000 406.350000 808.500000 407.650000 ;
      RECT 766.500000 406.350000 799.500000 407.650000 ;
      RECT 757.500000 406.350000 758.500000 407.650000 ;
      RECT 716.500000 406.350000 749.500000 407.650000 ;
      RECT 707.500000 406.350000 708.500000 407.650000 ;
      RECT 666.500000 406.350000 699.500000 407.650000 ;
      RECT 657.500000 406.350000 658.500000 407.650000 ;
      RECT 616.500000 406.350000 649.500000 407.650000 ;
      RECT 607.500000 406.350000 608.500000 407.650000 ;
      RECT 566.500000 406.350000 599.500000 407.650000 ;
      RECT 557.500000 406.350000 558.500000 407.650000 ;
      RECT 516.500000 406.350000 549.500000 407.650000 ;
      RECT 507.500000 406.350000 508.500000 407.650000 ;
      RECT 416.500000 406.350000 499.500000 407.650000 ;
      RECT 407.500000 406.350000 408.500000 407.650000 ;
      RECT 366.500000 406.350000 399.500000 407.650000 ;
      RECT 357.500000 406.350000 358.500000 407.650000 ;
      RECT 316.500000 406.350000 349.500000 407.650000 ;
      RECT 307.500000 406.350000 308.500000 407.650000 ;
      RECT 216.500000 406.350000 299.500000 407.650000 ;
      RECT 207.500000 406.350000 208.500000 407.650000 ;
      RECT 116.500000 406.350000 199.500000 407.650000 ;
      RECT 107.500000 406.350000 108.500000 407.650000 ;
      RECT 66.500000 406.350000 99.500000 407.650000 ;
      RECT 57.500000 406.350000 58.500000 407.650000 ;
      RECT 29.500000 406.350000 49.500000 407.650000 ;
      RECT 15.500000 406.350000 16.500000 407.650000 ;
      RECT 1157.500000 405.650000 1170.500000 406.350000 ;
      RECT 1107.500000 405.650000 1149.500000 406.350000 ;
      RECT 1057.500000 405.650000 1099.500000 406.350000 ;
      RECT 1007.500000 405.650000 1049.500000 406.350000 ;
      RECT 957.500000 405.650000 999.500000 406.350000 ;
      RECT 907.500000 405.650000 949.500000 406.350000 ;
      RECT 857.500000 405.650000 899.500000 406.350000 ;
      RECT 807.500000 405.650000 849.500000 406.350000 ;
      RECT 757.500000 405.650000 799.500000 406.350000 ;
      RECT 707.500000 405.650000 749.500000 406.350000 ;
      RECT 657.500000 405.650000 699.500000 406.350000 ;
      RECT 607.500000 405.650000 649.500000 406.350000 ;
      RECT 557.500000 405.650000 599.500000 406.350000 ;
      RECT 507.500000 405.650000 549.500000 406.350000 ;
      RECT 407.500000 405.650000 499.500000 406.350000 ;
      RECT 357.500000 405.650000 399.500000 406.350000 ;
      RECT 307.500000 405.650000 349.500000 406.350000 ;
      RECT 207.500000 405.650000 299.500000 406.350000 ;
      RECT 107.500000 405.650000 199.500000 406.350000 ;
      RECT 57.500000 405.650000 99.500000 406.350000 ;
      RECT 15.500000 405.650000 49.500000 406.350000 ;
      RECT 1183.500000 404.350000 1186.000000 407.650000 ;
      RECT 1169.500000 404.350000 1170.500000 405.650000 ;
      RECT 1116.500000 404.350000 1149.500000 405.650000 ;
      RECT 1107.500000 404.350000 1108.500000 405.650000 ;
      RECT 1066.500000 404.350000 1099.500000 405.650000 ;
      RECT 1057.500000 404.350000 1058.500000 405.650000 ;
      RECT 1016.500000 404.350000 1049.500000 405.650000 ;
      RECT 1007.500000 404.350000 1008.500000 405.650000 ;
      RECT 966.500000 404.350000 999.500000 405.650000 ;
      RECT 957.500000 404.350000 958.500000 405.650000 ;
      RECT 916.500000 404.350000 949.500000 405.650000 ;
      RECT 907.500000 404.350000 908.500000 405.650000 ;
      RECT 866.500000 404.350000 899.500000 405.650000 ;
      RECT 857.500000 404.350000 858.500000 405.650000 ;
      RECT 816.500000 404.350000 849.500000 405.650000 ;
      RECT 807.500000 404.350000 808.500000 405.650000 ;
      RECT 766.500000 404.350000 799.500000 405.650000 ;
      RECT 757.500000 404.350000 758.500000 405.650000 ;
      RECT 716.500000 404.350000 749.500000 405.650000 ;
      RECT 707.500000 404.350000 708.500000 405.650000 ;
      RECT 666.500000 404.350000 699.500000 405.650000 ;
      RECT 657.500000 404.350000 658.500000 405.650000 ;
      RECT 616.500000 404.350000 649.500000 405.650000 ;
      RECT 607.500000 404.350000 608.500000 405.650000 ;
      RECT 566.500000 404.350000 599.500000 405.650000 ;
      RECT 557.500000 404.350000 558.500000 405.650000 ;
      RECT 516.500000 404.350000 549.500000 405.650000 ;
      RECT 507.500000 404.350000 508.500000 405.650000 ;
      RECT 416.500000 404.350000 499.500000 405.650000 ;
      RECT 407.500000 404.350000 408.500000 405.650000 ;
      RECT 366.500000 404.350000 399.500000 405.650000 ;
      RECT 357.500000 404.350000 358.500000 405.650000 ;
      RECT 316.500000 404.350000 349.500000 405.650000 ;
      RECT 307.500000 404.350000 308.500000 405.650000 ;
      RECT 216.500000 404.350000 299.500000 405.650000 ;
      RECT 207.500000 404.350000 208.500000 405.650000 ;
      RECT 116.500000 404.350000 199.500000 405.650000 ;
      RECT 107.500000 404.350000 108.500000 405.650000 ;
      RECT 66.500000 404.350000 99.500000 405.650000 ;
      RECT 57.500000 404.350000 58.500000 405.650000 ;
      RECT 29.500000 404.350000 49.500000 405.650000 ;
      RECT 15.500000 404.350000 16.500000 405.650000 ;
      RECT 0.000000 404.350000 2.500000 407.650000 ;
      RECT 416.500000 403.730000 508.500000 404.350000 ;
      RECT 1169.500000 403.650000 1186.000000 404.350000 ;
      RECT 1116.500000 403.650000 1156.500000 404.350000 ;
      RECT 1066.500000 403.650000 1108.500000 404.350000 ;
      RECT 1016.500000 403.650000 1058.500000 404.350000 ;
      RECT 966.500000 403.650000 1008.500000 404.350000 ;
      RECT 916.500000 403.650000 958.500000 404.350000 ;
      RECT 866.500000 403.650000 908.500000 404.350000 ;
      RECT 816.500000 403.650000 858.500000 404.350000 ;
      RECT 766.500000 403.650000 808.500000 404.350000 ;
      RECT 716.500000 403.650000 758.500000 404.350000 ;
      RECT 666.500000 403.650000 708.500000 404.350000 ;
      RECT 616.500000 403.650000 658.500000 404.350000 ;
      RECT 566.500000 403.650000 608.500000 404.350000 ;
      RECT 516.500000 403.650000 558.500000 404.350000 ;
      RECT 466.500000 403.650000 508.500000 403.730000 ;
      RECT 366.500000 403.650000 408.500000 404.350000 ;
      RECT 316.500000 403.650000 358.500000 404.350000 ;
      RECT 216.500000 403.650000 308.500000 404.350000 ;
      RECT 116.500000 403.650000 208.500000 404.350000 ;
      RECT 66.500000 403.650000 108.500000 404.350000 ;
      RECT 29.500000 403.650000 58.500000 404.350000 ;
      RECT 0.000000 403.650000 16.500000 404.350000 ;
      RECT 1169.500000 402.350000 1170.500000 403.650000 ;
      RECT 1116.500000 402.350000 1149.500000 403.650000 ;
      RECT 1107.500000 402.350000 1108.500000 403.650000 ;
      RECT 1066.500000 402.350000 1099.500000 403.650000 ;
      RECT 1057.500000 402.350000 1058.500000 403.650000 ;
      RECT 1016.500000 402.350000 1049.500000 403.650000 ;
      RECT 1007.500000 402.350000 1008.500000 403.650000 ;
      RECT 966.500000 402.350000 999.500000 403.650000 ;
      RECT 957.500000 402.350000 958.500000 403.650000 ;
      RECT 916.500000 402.350000 949.500000 403.650000 ;
      RECT 907.500000 402.350000 908.500000 403.650000 ;
      RECT 866.500000 402.350000 899.500000 403.650000 ;
      RECT 857.500000 402.350000 858.500000 403.650000 ;
      RECT 816.500000 402.350000 849.500000 403.650000 ;
      RECT 807.500000 402.350000 808.500000 403.650000 ;
      RECT 766.500000 402.350000 799.500000 403.650000 ;
      RECT 757.500000 402.350000 758.500000 403.650000 ;
      RECT 716.500000 402.350000 749.500000 403.650000 ;
      RECT 707.500000 402.350000 708.500000 403.650000 ;
      RECT 666.500000 402.350000 699.500000 403.650000 ;
      RECT 657.500000 402.350000 658.500000 403.650000 ;
      RECT 616.500000 402.350000 649.500000 403.650000 ;
      RECT 607.500000 402.350000 608.500000 403.650000 ;
      RECT 566.500000 402.350000 599.500000 403.650000 ;
      RECT 557.500000 402.350000 558.500000 403.650000 ;
      RECT 516.500000 402.350000 549.500000 403.650000 ;
      RECT 507.500000 402.350000 508.500000 403.650000 ;
      RECT 416.500000 402.350000 458.500000 403.730000 ;
      RECT 407.500000 402.350000 408.500000 403.650000 ;
      RECT 366.500000 402.350000 399.500000 403.650000 ;
      RECT 357.500000 402.350000 358.500000 403.650000 ;
      RECT 316.500000 402.350000 349.500000 403.650000 ;
      RECT 307.500000 402.350000 308.500000 403.650000 ;
      RECT 216.500000 402.350000 249.500000 403.650000 ;
      RECT 207.500000 402.350000 208.500000 403.650000 ;
      RECT 116.500000 402.350000 149.500000 403.650000 ;
      RECT 107.500000 402.350000 108.500000 403.650000 ;
      RECT 66.500000 402.350000 99.500000 403.650000 ;
      RECT 57.500000 402.350000 58.500000 403.650000 ;
      RECT 29.500000 402.350000 49.500000 403.650000 ;
      RECT 15.500000 402.350000 16.500000 403.650000 ;
      RECT 1157.500000 401.650000 1170.500000 402.350000 ;
      RECT 1107.500000 401.650000 1149.500000 402.350000 ;
      RECT 1057.500000 401.650000 1099.500000 402.350000 ;
      RECT 1007.500000 401.650000 1049.500000 402.350000 ;
      RECT 957.500000 401.650000 999.500000 402.350000 ;
      RECT 907.500000 401.650000 949.500000 402.350000 ;
      RECT 857.500000 401.650000 899.500000 402.350000 ;
      RECT 807.500000 401.650000 849.500000 402.350000 ;
      RECT 757.500000 401.650000 799.500000 402.350000 ;
      RECT 707.500000 401.650000 749.500000 402.350000 ;
      RECT 657.500000 401.650000 699.500000 402.350000 ;
      RECT 607.500000 401.650000 649.500000 402.350000 ;
      RECT 557.500000 401.650000 599.500000 402.350000 ;
      RECT 507.500000 401.650000 549.500000 402.350000 ;
      RECT 407.500000 401.650000 458.500000 402.350000 ;
      RECT 357.500000 401.650000 399.500000 402.350000 ;
      RECT 307.500000 401.650000 349.500000 402.350000 ;
      RECT 257.500000 401.650000 299.500000 403.650000 ;
      RECT 207.500000 401.650000 249.500000 402.350000 ;
      RECT 157.500000 401.650000 199.500000 403.650000 ;
      RECT 107.500000 401.650000 149.500000 402.350000 ;
      RECT 57.500000 401.650000 99.500000 402.350000 ;
      RECT 15.500000 401.650000 49.500000 402.350000 ;
      RECT 1183.500000 400.350000 1186.000000 403.650000 ;
      RECT 1169.500000 400.350000 1170.500000 401.650000 ;
      RECT 1116.500000 400.350000 1149.500000 401.650000 ;
      RECT 1107.500000 400.350000 1108.500000 401.650000 ;
      RECT 1066.500000 400.350000 1099.500000 401.650000 ;
      RECT 1057.500000 400.350000 1058.500000 401.650000 ;
      RECT 1016.500000 400.350000 1049.500000 401.650000 ;
      RECT 1007.500000 400.350000 1008.500000 401.650000 ;
      RECT 966.500000 400.350000 999.500000 401.650000 ;
      RECT 957.500000 400.350000 958.500000 401.650000 ;
      RECT 916.500000 400.350000 949.500000 401.650000 ;
      RECT 907.500000 400.350000 908.500000 401.650000 ;
      RECT 866.500000 400.350000 899.500000 401.650000 ;
      RECT 857.500000 400.350000 858.500000 401.650000 ;
      RECT 816.500000 400.350000 849.500000 401.650000 ;
      RECT 807.500000 400.350000 808.500000 401.650000 ;
      RECT 766.500000 400.350000 799.500000 401.650000 ;
      RECT 757.500000 400.350000 758.500000 401.650000 ;
      RECT 716.500000 400.350000 749.500000 401.650000 ;
      RECT 707.500000 400.350000 708.500000 401.650000 ;
      RECT 666.500000 400.350000 699.500000 401.650000 ;
      RECT 657.500000 400.350000 658.500000 401.650000 ;
      RECT 616.500000 400.350000 649.500000 401.650000 ;
      RECT 607.500000 400.350000 608.500000 401.650000 ;
      RECT 566.500000 400.350000 599.500000 401.650000 ;
      RECT 557.500000 400.350000 558.500000 401.650000 ;
      RECT 516.500000 400.350000 549.500000 401.650000 ;
      RECT 507.500000 400.350000 508.500000 401.650000 ;
      RECT 466.500000 400.350000 499.500000 403.650000 ;
      RECT 407.500000 400.350000 408.500000 401.650000 ;
      RECT 366.500000 400.350000 399.500000 401.650000 ;
      RECT 357.500000 400.350000 358.500000 401.650000 ;
      RECT 316.500000 400.350000 349.500000 401.650000 ;
      RECT 307.500000 400.350000 308.500000 401.650000 ;
      RECT 266.500000 400.350000 299.500000 401.650000 ;
      RECT 257.500000 400.350000 258.500000 401.650000 ;
      RECT 216.500000 400.350000 249.500000 401.650000 ;
      RECT 207.500000 400.350000 208.500000 401.650000 ;
      RECT 166.500000 400.350000 199.500000 401.650000 ;
      RECT 157.500000 400.350000 158.500000 401.650000 ;
      RECT 116.500000 400.350000 149.500000 401.650000 ;
      RECT 107.500000 400.350000 108.500000 401.650000 ;
      RECT 66.500000 400.350000 99.500000 401.650000 ;
      RECT 57.500000 400.350000 58.500000 401.650000 ;
      RECT 29.500000 400.350000 49.500000 401.650000 ;
      RECT 15.500000 400.350000 16.500000 401.650000 ;
      RECT 0.000000 400.350000 2.500000 403.650000 ;
      RECT 466.500000 399.730000 508.500000 400.350000 ;
      RECT 416.500000 399.730000 458.500000 401.650000 ;
      RECT 1169.500000 399.650000 1186.000000 400.350000 ;
      RECT 1116.500000 399.650000 1156.500000 400.350000 ;
      RECT 1066.500000 399.650000 1108.500000 400.350000 ;
      RECT 1016.500000 399.650000 1058.500000 400.350000 ;
      RECT 966.500000 399.650000 1008.500000 400.350000 ;
      RECT 916.500000 399.650000 958.500000 400.350000 ;
      RECT 866.500000 399.650000 908.500000 400.350000 ;
      RECT 816.500000 399.650000 858.500000 400.350000 ;
      RECT 766.500000 399.650000 808.500000 400.350000 ;
      RECT 716.500000 399.650000 758.500000 400.350000 ;
      RECT 666.500000 399.650000 708.500000 400.350000 ;
      RECT 616.500000 399.650000 658.500000 400.350000 ;
      RECT 566.500000 399.650000 608.500000 400.350000 ;
      RECT 516.500000 399.650000 558.500000 400.350000 ;
      RECT 416.500000 399.650000 508.500000 399.730000 ;
      RECT 366.500000 399.650000 408.500000 400.350000 ;
      RECT 316.500000 399.650000 358.500000 400.350000 ;
      RECT 266.500000 399.650000 308.500000 400.350000 ;
      RECT 216.500000 399.650000 258.500000 400.350000 ;
      RECT 166.500000 399.650000 208.500000 400.350000 ;
      RECT 116.500000 399.650000 158.500000 400.350000 ;
      RECT 66.500000 399.650000 108.500000 400.350000 ;
      RECT 29.500000 399.650000 58.500000 400.350000 ;
      RECT 0.000000 399.650000 16.500000 400.350000 ;
      RECT 1169.500000 398.350000 1170.500000 399.650000 ;
      RECT 1116.500000 398.350000 1149.500000 399.650000 ;
      RECT 1107.500000 398.350000 1108.500000 399.650000 ;
      RECT 1066.500000 398.350000 1099.500000 399.650000 ;
      RECT 1057.500000 398.350000 1058.500000 399.650000 ;
      RECT 1016.500000 398.350000 1049.500000 399.650000 ;
      RECT 1007.500000 398.350000 1008.500000 399.650000 ;
      RECT 966.500000 398.350000 999.500000 399.650000 ;
      RECT 957.500000 398.350000 958.500000 399.650000 ;
      RECT 916.500000 398.350000 949.500000 399.650000 ;
      RECT 907.500000 398.350000 908.500000 399.650000 ;
      RECT 866.500000 398.350000 899.500000 399.650000 ;
      RECT 857.500000 398.350000 858.500000 399.650000 ;
      RECT 816.500000 398.350000 849.500000 399.650000 ;
      RECT 807.500000 398.350000 808.500000 399.650000 ;
      RECT 766.500000 398.350000 799.500000 399.650000 ;
      RECT 757.500000 398.350000 758.500000 399.650000 ;
      RECT 716.500000 398.350000 749.500000 399.650000 ;
      RECT 707.500000 398.350000 708.500000 399.650000 ;
      RECT 666.500000 398.350000 699.500000 399.650000 ;
      RECT 657.500000 398.350000 658.500000 399.650000 ;
      RECT 616.500000 398.350000 649.500000 399.650000 ;
      RECT 607.500000 398.350000 608.500000 399.650000 ;
      RECT 566.500000 398.350000 599.500000 399.650000 ;
      RECT 557.500000 398.350000 558.500000 399.650000 ;
      RECT 516.500000 398.350000 549.500000 399.650000 ;
      RECT 507.500000 398.350000 508.500000 399.650000 ;
      RECT 416.500000 398.350000 449.500000 399.650000 ;
      RECT 407.500000 398.350000 408.500000 399.650000 ;
      RECT 366.500000 398.350000 399.500000 399.650000 ;
      RECT 357.500000 398.350000 358.500000 399.650000 ;
      RECT 316.500000 398.350000 349.500000 399.650000 ;
      RECT 307.500000 398.350000 308.500000 399.650000 ;
      RECT 266.500000 398.350000 299.500000 399.650000 ;
      RECT 257.500000 398.350000 258.500000 399.650000 ;
      RECT 216.500000 398.350000 249.500000 399.650000 ;
      RECT 207.500000 398.350000 208.500000 399.650000 ;
      RECT 166.500000 398.350000 199.500000 399.650000 ;
      RECT 157.500000 398.350000 158.500000 399.650000 ;
      RECT 116.500000 398.350000 149.500000 399.650000 ;
      RECT 107.500000 398.350000 108.500000 399.650000 ;
      RECT 66.500000 398.350000 99.500000 399.650000 ;
      RECT 57.500000 398.350000 58.500000 399.650000 ;
      RECT 29.500000 398.350000 49.500000 399.650000 ;
      RECT 15.500000 398.350000 16.500000 399.650000 ;
      RECT 1157.500000 397.650000 1170.500000 398.350000 ;
      RECT 1107.500000 397.650000 1149.500000 398.350000 ;
      RECT 1057.500000 397.650000 1099.500000 398.350000 ;
      RECT 1007.500000 397.650000 1049.500000 398.350000 ;
      RECT 957.500000 397.650000 999.500000 398.350000 ;
      RECT 907.500000 397.650000 949.500000 398.350000 ;
      RECT 857.500000 397.650000 899.500000 398.350000 ;
      RECT 807.500000 397.650000 849.500000 398.350000 ;
      RECT 757.500000 397.650000 799.500000 398.350000 ;
      RECT 707.500000 397.650000 749.500000 398.350000 ;
      RECT 657.500000 397.650000 699.500000 398.350000 ;
      RECT 607.500000 397.650000 649.500000 398.350000 ;
      RECT 557.500000 397.650000 599.500000 398.350000 ;
      RECT 507.500000 397.650000 549.500000 398.350000 ;
      RECT 457.500000 397.650000 499.500000 399.650000 ;
      RECT 407.500000 397.650000 449.500000 398.350000 ;
      RECT 357.500000 397.650000 399.500000 398.350000 ;
      RECT 307.500000 397.650000 349.500000 398.350000 ;
      RECT 257.500000 397.650000 299.500000 398.350000 ;
      RECT 207.500000 397.650000 249.500000 398.350000 ;
      RECT 157.500000 397.650000 199.500000 398.350000 ;
      RECT 107.500000 397.650000 149.500000 398.350000 ;
      RECT 57.500000 397.650000 99.500000 398.350000 ;
      RECT 15.500000 397.650000 49.500000 398.350000 ;
      RECT 1183.500000 396.350000 1186.000000 399.650000 ;
      RECT 1169.500000 396.350000 1170.500000 397.650000 ;
      RECT 1116.500000 396.350000 1149.500000 397.650000 ;
      RECT 1107.500000 396.350000 1108.500000 397.650000 ;
      RECT 1066.500000 396.350000 1099.500000 397.650000 ;
      RECT 1057.500000 396.350000 1058.500000 397.650000 ;
      RECT 1016.500000 396.350000 1049.500000 397.650000 ;
      RECT 1007.500000 396.350000 1008.500000 397.650000 ;
      RECT 966.500000 396.350000 999.500000 397.650000 ;
      RECT 957.500000 396.350000 958.500000 397.650000 ;
      RECT 916.500000 396.350000 949.500000 397.650000 ;
      RECT 907.500000 396.350000 908.500000 397.650000 ;
      RECT 866.500000 396.350000 899.500000 397.650000 ;
      RECT 857.500000 396.350000 858.500000 397.650000 ;
      RECT 816.500000 396.350000 849.500000 397.650000 ;
      RECT 807.500000 396.350000 808.500000 397.650000 ;
      RECT 766.500000 396.350000 799.500000 397.650000 ;
      RECT 757.500000 396.350000 758.500000 397.650000 ;
      RECT 716.500000 396.350000 749.500000 397.650000 ;
      RECT 707.500000 396.350000 708.500000 397.650000 ;
      RECT 666.500000 396.350000 699.500000 397.650000 ;
      RECT 657.500000 396.350000 658.500000 397.650000 ;
      RECT 616.500000 396.350000 649.500000 397.650000 ;
      RECT 607.500000 396.350000 608.500000 397.650000 ;
      RECT 566.500000 396.350000 599.500000 397.650000 ;
      RECT 557.500000 396.350000 558.500000 397.650000 ;
      RECT 516.500000 396.350000 549.500000 397.650000 ;
      RECT 507.500000 396.350000 508.500000 397.650000 ;
      RECT 466.500000 396.350000 499.500000 397.650000 ;
      RECT 457.500000 396.350000 458.500000 397.650000 ;
      RECT 416.500000 396.350000 449.500000 397.650000 ;
      RECT 407.500000 396.350000 408.500000 397.650000 ;
      RECT 366.500000 396.350000 399.500000 397.650000 ;
      RECT 357.500000 396.350000 358.500000 397.650000 ;
      RECT 316.500000 396.350000 349.500000 397.650000 ;
      RECT 307.500000 396.350000 308.500000 397.650000 ;
      RECT 266.500000 396.350000 299.500000 397.650000 ;
      RECT 257.500000 396.350000 258.500000 397.650000 ;
      RECT 216.500000 396.350000 249.500000 397.650000 ;
      RECT 207.500000 396.350000 208.500000 397.650000 ;
      RECT 166.500000 396.350000 199.500000 397.650000 ;
      RECT 157.500000 396.350000 158.500000 397.650000 ;
      RECT 116.500000 396.350000 149.500000 397.650000 ;
      RECT 107.500000 396.350000 108.500000 397.650000 ;
      RECT 66.500000 396.350000 99.500000 397.650000 ;
      RECT 57.500000 396.350000 58.500000 397.650000 ;
      RECT 29.500000 396.350000 49.500000 397.650000 ;
      RECT 15.500000 396.350000 16.500000 397.650000 ;
      RECT 0.000000 396.350000 2.500000 399.650000 ;
      RECT 1169.500000 395.650000 1186.000000 396.350000 ;
      RECT 1116.500000 395.650000 1156.500000 396.350000 ;
      RECT 1066.500000 395.650000 1108.500000 396.350000 ;
      RECT 1016.500000 395.650000 1058.500000 396.350000 ;
      RECT 966.500000 395.650000 1008.500000 396.350000 ;
      RECT 916.500000 395.650000 958.500000 396.350000 ;
      RECT 866.500000 395.650000 908.500000 396.350000 ;
      RECT 816.500000 395.650000 858.500000 396.350000 ;
      RECT 766.500000 395.650000 808.500000 396.350000 ;
      RECT 716.500000 395.650000 758.500000 396.350000 ;
      RECT 666.500000 395.650000 708.500000 396.350000 ;
      RECT 616.500000 395.650000 658.500000 396.350000 ;
      RECT 566.500000 395.650000 608.500000 396.350000 ;
      RECT 516.500000 395.650000 558.500000 396.350000 ;
      RECT 466.500000 395.650000 508.500000 396.350000 ;
      RECT 416.500000 395.650000 458.500000 396.350000 ;
      RECT 366.500000 395.650000 408.500000 396.350000 ;
      RECT 316.500000 395.650000 358.500000 396.350000 ;
      RECT 266.500000 395.650000 308.500000 396.350000 ;
      RECT 216.500000 395.650000 258.500000 396.350000 ;
      RECT 166.500000 395.650000 208.500000 396.350000 ;
      RECT 116.500000 395.650000 158.500000 396.350000 ;
      RECT 66.500000 395.650000 108.500000 396.350000 ;
      RECT 29.500000 395.650000 58.500000 396.350000 ;
      RECT 0.000000 395.650000 16.500000 396.350000 ;
      RECT 1169.500000 394.350000 1170.500000 395.650000 ;
      RECT 1116.500000 394.350000 1149.500000 395.650000 ;
      RECT 1107.500000 394.350000 1108.500000 395.650000 ;
      RECT 1066.500000 394.350000 1099.500000 395.650000 ;
      RECT 1057.500000 394.350000 1058.500000 395.650000 ;
      RECT 1016.500000 394.350000 1049.500000 395.650000 ;
      RECT 1007.500000 394.350000 1008.500000 395.650000 ;
      RECT 966.500000 394.350000 999.500000 395.650000 ;
      RECT 957.500000 394.350000 958.500000 395.650000 ;
      RECT 916.500000 394.350000 949.500000 395.650000 ;
      RECT 907.500000 394.350000 908.500000 395.650000 ;
      RECT 866.500000 394.350000 899.500000 395.650000 ;
      RECT 857.500000 394.350000 858.500000 395.650000 ;
      RECT 816.500000 394.350000 849.500000 395.650000 ;
      RECT 807.500000 394.350000 808.500000 395.650000 ;
      RECT 766.500000 394.350000 799.500000 395.650000 ;
      RECT 757.500000 394.350000 758.500000 395.650000 ;
      RECT 716.500000 394.350000 749.500000 395.650000 ;
      RECT 707.500000 394.350000 708.500000 395.650000 ;
      RECT 666.500000 394.350000 699.500000 395.650000 ;
      RECT 657.500000 394.350000 658.500000 395.650000 ;
      RECT 616.500000 394.350000 649.500000 395.650000 ;
      RECT 607.500000 394.350000 608.500000 395.650000 ;
      RECT 566.500000 394.350000 599.500000 395.650000 ;
      RECT 557.500000 394.350000 558.500000 395.650000 ;
      RECT 516.500000 394.350000 549.500000 395.650000 ;
      RECT 507.500000 394.350000 508.500000 395.650000 ;
      RECT 466.500000 394.350000 499.500000 395.650000 ;
      RECT 457.500000 394.350000 458.500000 395.650000 ;
      RECT 416.500000 394.350000 449.500000 395.650000 ;
      RECT 407.500000 394.350000 408.500000 395.650000 ;
      RECT 366.500000 394.350000 399.500000 395.650000 ;
      RECT 357.500000 394.350000 358.500000 395.650000 ;
      RECT 316.500000 394.350000 349.500000 395.650000 ;
      RECT 307.500000 394.350000 308.500000 395.650000 ;
      RECT 266.500000 394.350000 299.500000 395.650000 ;
      RECT 257.500000 394.350000 258.500000 395.650000 ;
      RECT 216.500000 394.350000 249.500000 395.650000 ;
      RECT 207.500000 394.350000 208.500000 395.650000 ;
      RECT 166.500000 394.350000 199.500000 395.650000 ;
      RECT 157.500000 394.350000 158.500000 395.650000 ;
      RECT 116.500000 394.350000 149.500000 395.650000 ;
      RECT 107.500000 394.350000 108.500000 395.650000 ;
      RECT 66.500000 394.350000 99.500000 395.650000 ;
      RECT 57.500000 394.350000 58.500000 395.650000 ;
      RECT 29.500000 394.350000 49.500000 395.650000 ;
      RECT 15.500000 394.350000 16.500000 395.650000 ;
      RECT 1157.500000 393.650000 1170.500000 394.350000 ;
      RECT 1107.500000 393.650000 1149.500000 394.350000 ;
      RECT 1057.500000 393.650000 1099.500000 394.350000 ;
      RECT 1007.500000 393.650000 1049.500000 394.350000 ;
      RECT 957.500000 393.650000 999.500000 394.350000 ;
      RECT 907.500000 393.650000 949.500000 394.350000 ;
      RECT 857.500000 393.650000 899.500000 394.350000 ;
      RECT 807.500000 393.650000 849.500000 394.350000 ;
      RECT 757.500000 393.650000 799.500000 394.350000 ;
      RECT 707.500000 393.650000 749.500000 394.350000 ;
      RECT 657.500000 393.650000 699.500000 394.350000 ;
      RECT 607.500000 393.650000 649.500000 394.350000 ;
      RECT 557.500000 393.650000 599.500000 394.350000 ;
      RECT 507.500000 393.650000 549.500000 394.350000 ;
      RECT 457.500000 393.650000 499.500000 394.350000 ;
      RECT 407.500000 393.650000 449.500000 394.350000 ;
      RECT 357.500000 393.650000 399.500000 394.350000 ;
      RECT 307.500000 393.650000 349.500000 394.350000 ;
      RECT 257.500000 393.650000 299.500000 394.350000 ;
      RECT 207.500000 393.650000 249.500000 394.350000 ;
      RECT 157.500000 393.650000 199.500000 394.350000 ;
      RECT 107.500000 393.650000 149.500000 394.350000 ;
      RECT 57.500000 393.650000 99.500000 394.350000 ;
      RECT 15.500000 393.650000 49.500000 394.350000 ;
      RECT 1183.500000 392.350000 1186.000000 395.650000 ;
      RECT 1169.500000 392.350000 1170.500000 393.650000 ;
      RECT 1116.500000 392.350000 1149.500000 393.650000 ;
      RECT 1107.500000 392.350000 1108.500000 393.650000 ;
      RECT 1066.500000 392.350000 1099.500000 393.650000 ;
      RECT 1057.500000 392.350000 1058.500000 393.650000 ;
      RECT 1016.500000 392.350000 1049.500000 393.650000 ;
      RECT 1007.500000 392.350000 1008.500000 393.650000 ;
      RECT 966.500000 392.350000 999.500000 393.650000 ;
      RECT 957.500000 392.350000 958.500000 393.650000 ;
      RECT 916.500000 392.350000 949.500000 393.650000 ;
      RECT 907.500000 392.350000 908.500000 393.650000 ;
      RECT 866.500000 392.350000 899.500000 393.650000 ;
      RECT 857.500000 392.350000 858.500000 393.650000 ;
      RECT 816.500000 392.350000 849.500000 393.650000 ;
      RECT 807.500000 392.350000 808.500000 393.650000 ;
      RECT 766.500000 392.350000 799.500000 393.650000 ;
      RECT 757.500000 392.350000 758.500000 393.650000 ;
      RECT 716.500000 392.350000 749.500000 393.650000 ;
      RECT 707.500000 392.350000 708.500000 393.650000 ;
      RECT 666.500000 392.350000 699.500000 393.650000 ;
      RECT 657.500000 392.350000 658.500000 393.650000 ;
      RECT 616.500000 392.350000 649.500000 393.650000 ;
      RECT 607.500000 392.350000 608.500000 393.650000 ;
      RECT 566.500000 392.350000 599.500000 393.650000 ;
      RECT 557.500000 392.350000 558.500000 393.650000 ;
      RECT 516.500000 392.350000 549.500000 393.650000 ;
      RECT 507.500000 392.350000 508.500000 393.650000 ;
      RECT 466.500000 392.350000 499.500000 393.650000 ;
      RECT 457.500000 392.350000 458.500000 393.650000 ;
      RECT 416.500000 392.350000 449.500000 393.650000 ;
      RECT 407.500000 392.350000 408.500000 393.650000 ;
      RECT 366.500000 392.350000 399.500000 393.650000 ;
      RECT 357.500000 392.350000 358.500000 393.650000 ;
      RECT 316.500000 392.350000 349.500000 393.650000 ;
      RECT 307.500000 392.350000 308.500000 393.650000 ;
      RECT 266.500000 392.350000 299.500000 393.650000 ;
      RECT 257.500000 392.350000 258.500000 393.650000 ;
      RECT 216.500000 392.350000 249.500000 393.650000 ;
      RECT 207.500000 392.350000 208.500000 393.650000 ;
      RECT 166.500000 392.350000 199.500000 393.650000 ;
      RECT 157.500000 392.350000 158.500000 393.650000 ;
      RECT 116.500000 392.350000 149.500000 393.650000 ;
      RECT 107.500000 392.350000 108.500000 393.650000 ;
      RECT 66.500000 392.350000 99.500000 393.650000 ;
      RECT 57.500000 392.350000 58.500000 393.650000 ;
      RECT 29.500000 392.350000 49.500000 393.650000 ;
      RECT 15.500000 392.350000 16.500000 393.650000 ;
      RECT 0.000000 392.350000 2.500000 395.650000 ;
      RECT 1169.500000 391.650000 1186.000000 392.350000 ;
      RECT 1116.500000 391.650000 1156.500000 392.350000 ;
      RECT 1066.500000 391.650000 1108.500000 392.350000 ;
      RECT 1016.500000 391.650000 1058.500000 392.350000 ;
      RECT 966.500000 391.650000 1008.500000 392.350000 ;
      RECT 916.500000 391.650000 958.500000 392.350000 ;
      RECT 866.500000 391.650000 908.500000 392.350000 ;
      RECT 816.500000 391.650000 858.500000 392.350000 ;
      RECT 766.500000 391.650000 808.500000 392.350000 ;
      RECT 716.500000 391.650000 758.500000 392.350000 ;
      RECT 666.500000 391.650000 708.500000 392.350000 ;
      RECT 616.500000 391.650000 658.500000 392.350000 ;
      RECT 566.500000 391.650000 608.500000 392.350000 ;
      RECT 516.500000 391.650000 558.500000 392.350000 ;
      RECT 466.500000 391.650000 508.500000 392.350000 ;
      RECT 416.500000 391.650000 458.500000 392.350000 ;
      RECT 366.500000 391.650000 408.500000 392.350000 ;
      RECT 316.500000 391.650000 358.500000 392.350000 ;
      RECT 266.500000 391.650000 308.500000 392.350000 ;
      RECT 216.500000 391.650000 258.500000 392.350000 ;
      RECT 166.500000 391.650000 208.500000 392.350000 ;
      RECT 116.500000 391.650000 158.500000 392.350000 ;
      RECT 66.500000 391.650000 108.500000 392.350000 ;
      RECT 29.500000 391.650000 58.500000 392.350000 ;
      RECT 0.000000 391.650000 16.500000 392.350000 ;
      RECT 1169.500000 390.350000 1170.500000 391.650000 ;
      RECT 1116.500000 390.350000 1149.500000 391.650000 ;
      RECT 1107.500000 390.350000 1108.500000 391.650000 ;
      RECT 1066.500000 390.350000 1099.500000 391.650000 ;
      RECT 1057.500000 390.350000 1058.500000 391.650000 ;
      RECT 1016.500000 390.350000 1049.500000 391.650000 ;
      RECT 1007.500000 390.350000 1008.500000 391.650000 ;
      RECT 966.500000 390.350000 999.500000 391.650000 ;
      RECT 957.500000 390.350000 958.500000 391.650000 ;
      RECT 916.500000 390.350000 949.500000 391.650000 ;
      RECT 907.500000 390.350000 908.500000 391.650000 ;
      RECT 866.500000 390.350000 899.500000 391.650000 ;
      RECT 857.500000 390.350000 858.500000 391.650000 ;
      RECT 816.500000 390.350000 849.500000 391.650000 ;
      RECT 807.500000 390.350000 808.500000 391.650000 ;
      RECT 766.500000 390.350000 799.500000 391.650000 ;
      RECT 757.500000 390.350000 758.500000 391.650000 ;
      RECT 716.500000 390.350000 749.500000 391.650000 ;
      RECT 707.500000 390.350000 708.500000 391.650000 ;
      RECT 666.500000 390.350000 699.500000 391.650000 ;
      RECT 657.500000 390.350000 658.500000 391.650000 ;
      RECT 616.500000 390.350000 649.500000 391.650000 ;
      RECT 607.500000 390.350000 608.500000 391.650000 ;
      RECT 566.500000 390.350000 599.500000 391.650000 ;
      RECT 557.500000 390.350000 558.500000 391.650000 ;
      RECT 516.500000 390.350000 549.500000 391.650000 ;
      RECT 507.500000 390.350000 508.500000 391.650000 ;
      RECT 466.500000 390.350000 499.500000 391.650000 ;
      RECT 457.500000 390.350000 458.500000 391.650000 ;
      RECT 416.500000 390.350000 449.500000 391.650000 ;
      RECT 407.500000 390.350000 408.500000 391.650000 ;
      RECT 366.500000 390.350000 399.500000 391.650000 ;
      RECT 357.500000 390.350000 358.500000 391.650000 ;
      RECT 316.500000 390.350000 349.500000 391.650000 ;
      RECT 307.500000 390.350000 308.500000 391.650000 ;
      RECT 266.500000 390.350000 299.500000 391.650000 ;
      RECT 257.500000 390.350000 258.500000 391.650000 ;
      RECT 216.500000 390.350000 249.500000 391.650000 ;
      RECT 207.500000 390.350000 208.500000 391.650000 ;
      RECT 166.500000 390.350000 199.500000 391.650000 ;
      RECT 157.500000 390.350000 158.500000 391.650000 ;
      RECT 116.500000 390.350000 149.500000 391.650000 ;
      RECT 107.500000 390.350000 108.500000 391.650000 ;
      RECT 66.500000 390.350000 99.500000 391.650000 ;
      RECT 57.500000 390.350000 58.500000 391.650000 ;
      RECT 29.500000 390.350000 49.500000 391.650000 ;
      RECT 15.500000 390.350000 16.500000 391.650000 ;
      RECT 1157.500000 389.650000 1170.500000 390.350000 ;
      RECT 1107.500000 389.650000 1149.500000 390.350000 ;
      RECT 1057.500000 389.650000 1099.500000 390.350000 ;
      RECT 1007.500000 389.650000 1049.500000 390.350000 ;
      RECT 957.500000 389.650000 999.500000 390.350000 ;
      RECT 907.500000 389.650000 949.500000 390.350000 ;
      RECT 857.500000 389.650000 899.500000 390.350000 ;
      RECT 807.500000 389.650000 849.500000 390.350000 ;
      RECT 757.500000 389.650000 799.500000 390.350000 ;
      RECT 707.500000 389.650000 749.500000 390.350000 ;
      RECT 657.500000 389.650000 699.500000 390.350000 ;
      RECT 607.500000 389.650000 649.500000 390.350000 ;
      RECT 557.500000 389.650000 599.500000 390.350000 ;
      RECT 507.500000 389.650000 549.500000 390.350000 ;
      RECT 457.500000 389.650000 499.500000 390.350000 ;
      RECT 407.500000 389.650000 449.500000 390.350000 ;
      RECT 357.500000 389.650000 399.500000 390.350000 ;
      RECT 307.500000 389.650000 349.500000 390.350000 ;
      RECT 257.500000 389.650000 299.500000 390.350000 ;
      RECT 207.500000 389.650000 249.500000 390.350000 ;
      RECT 157.500000 389.650000 199.500000 390.350000 ;
      RECT 107.500000 389.650000 149.500000 390.350000 ;
      RECT 57.500000 389.650000 99.500000 390.350000 ;
      RECT 15.500000 389.650000 49.500000 390.350000 ;
      RECT 1183.500000 388.350000 1186.000000 391.650000 ;
      RECT 1169.500000 388.350000 1170.500000 389.650000 ;
      RECT 1116.500000 388.350000 1149.500000 389.650000 ;
      RECT 1107.500000 388.350000 1108.500000 389.650000 ;
      RECT 1066.500000 388.350000 1099.500000 389.650000 ;
      RECT 1057.500000 388.350000 1058.500000 389.650000 ;
      RECT 1016.500000 388.350000 1049.500000 389.650000 ;
      RECT 1007.500000 388.350000 1008.500000 389.650000 ;
      RECT 966.500000 388.350000 999.500000 389.650000 ;
      RECT 957.500000 388.350000 958.500000 389.650000 ;
      RECT 916.500000 388.350000 949.500000 389.650000 ;
      RECT 907.500000 388.350000 908.500000 389.650000 ;
      RECT 866.500000 388.350000 899.500000 389.650000 ;
      RECT 857.500000 388.350000 858.500000 389.650000 ;
      RECT 816.500000 388.350000 849.500000 389.650000 ;
      RECT 807.500000 388.350000 808.500000 389.650000 ;
      RECT 766.500000 388.350000 799.500000 389.650000 ;
      RECT 757.500000 388.350000 758.500000 389.650000 ;
      RECT 716.500000 388.350000 749.500000 389.650000 ;
      RECT 707.500000 388.350000 708.500000 389.650000 ;
      RECT 666.500000 388.350000 699.500000 389.650000 ;
      RECT 657.500000 388.350000 658.500000 389.650000 ;
      RECT 616.500000 388.350000 649.500000 389.650000 ;
      RECT 607.500000 388.350000 608.500000 389.650000 ;
      RECT 566.500000 388.350000 599.500000 389.650000 ;
      RECT 557.500000 388.350000 558.500000 389.650000 ;
      RECT 516.500000 388.350000 549.500000 389.650000 ;
      RECT 507.500000 388.350000 508.500000 389.650000 ;
      RECT 466.500000 388.350000 499.500000 389.650000 ;
      RECT 457.500000 388.350000 458.500000 389.650000 ;
      RECT 416.500000 388.350000 449.500000 389.650000 ;
      RECT 407.500000 388.350000 408.500000 389.650000 ;
      RECT 366.500000 388.350000 399.500000 389.650000 ;
      RECT 357.500000 388.350000 358.500000 389.650000 ;
      RECT 316.500000 388.350000 349.500000 389.650000 ;
      RECT 307.500000 388.350000 308.500000 389.650000 ;
      RECT 266.500000 388.350000 299.500000 389.650000 ;
      RECT 257.500000 388.350000 258.500000 389.650000 ;
      RECT 216.500000 388.350000 249.500000 389.650000 ;
      RECT 207.500000 388.350000 208.500000 389.650000 ;
      RECT 166.500000 388.350000 199.500000 389.650000 ;
      RECT 157.500000 388.350000 158.500000 389.650000 ;
      RECT 116.500000 388.350000 149.500000 389.650000 ;
      RECT 107.500000 388.350000 108.500000 389.650000 ;
      RECT 66.500000 388.350000 99.500000 389.650000 ;
      RECT 57.500000 388.350000 58.500000 389.650000 ;
      RECT 29.500000 388.350000 49.500000 389.650000 ;
      RECT 15.500000 388.350000 16.500000 389.650000 ;
      RECT 0.000000 388.350000 2.500000 391.650000 ;
      RECT 1169.500000 387.650000 1186.000000 388.350000 ;
      RECT 1116.500000 387.650000 1156.500000 388.350000 ;
      RECT 1066.500000 387.650000 1108.500000 388.350000 ;
      RECT 1016.500000 387.650000 1058.500000 388.350000 ;
      RECT 966.500000 387.650000 1008.500000 388.350000 ;
      RECT 916.500000 387.650000 958.500000 388.350000 ;
      RECT 866.500000 387.650000 908.500000 388.350000 ;
      RECT 816.500000 387.650000 858.500000 388.350000 ;
      RECT 766.500000 387.650000 808.500000 388.350000 ;
      RECT 716.500000 387.650000 758.500000 388.350000 ;
      RECT 666.500000 387.650000 708.500000 388.350000 ;
      RECT 616.500000 387.650000 658.500000 388.350000 ;
      RECT 566.500000 387.650000 608.500000 388.350000 ;
      RECT 516.500000 387.650000 558.500000 388.350000 ;
      RECT 466.500000 387.650000 508.500000 388.350000 ;
      RECT 416.500000 387.650000 458.500000 388.350000 ;
      RECT 366.500000 387.650000 408.500000 388.350000 ;
      RECT 316.500000 387.650000 358.500000 388.350000 ;
      RECT 266.500000 387.650000 308.500000 388.350000 ;
      RECT 216.500000 387.650000 258.500000 388.350000 ;
      RECT 166.500000 387.650000 208.500000 388.350000 ;
      RECT 116.500000 387.650000 158.500000 388.350000 ;
      RECT 66.500000 387.650000 108.500000 388.350000 ;
      RECT 29.500000 387.650000 58.500000 388.350000 ;
      RECT 0.000000 387.650000 16.500000 388.350000 ;
      RECT 1169.500000 386.350000 1170.500000 387.650000 ;
      RECT 1116.500000 386.350000 1149.500000 387.650000 ;
      RECT 1107.500000 386.350000 1108.500000 387.650000 ;
      RECT 1066.500000 386.350000 1099.500000 387.650000 ;
      RECT 1057.500000 386.350000 1058.500000 387.650000 ;
      RECT 1016.500000 386.350000 1049.500000 387.650000 ;
      RECT 1007.500000 386.350000 1008.500000 387.650000 ;
      RECT 966.500000 386.350000 999.500000 387.650000 ;
      RECT 957.500000 386.350000 958.500000 387.650000 ;
      RECT 916.500000 386.350000 949.500000 387.650000 ;
      RECT 907.500000 386.350000 908.500000 387.650000 ;
      RECT 866.500000 386.350000 899.500000 387.650000 ;
      RECT 857.500000 386.350000 858.500000 387.650000 ;
      RECT 816.500000 386.350000 849.500000 387.650000 ;
      RECT 807.500000 386.350000 808.500000 387.650000 ;
      RECT 766.500000 386.350000 799.500000 387.650000 ;
      RECT 757.500000 386.350000 758.500000 387.650000 ;
      RECT 716.500000 386.350000 749.500000 387.650000 ;
      RECT 707.500000 386.350000 708.500000 387.650000 ;
      RECT 666.500000 386.350000 699.500000 387.650000 ;
      RECT 657.500000 386.350000 658.500000 387.650000 ;
      RECT 616.500000 386.350000 649.500000 387.650000 ;
      RECT 607.500000 386.350000 608.500000 387.650000 ;
      RECT 566.500000 386.350000 599.500000 387.650000 ;
      RECT 557.500000 386.350000 558.500000 387.650000 ;
      RECT 516.500000 386.350000 549.500000 387.650000 ;
      RECT 507.500000 386.350000 508.500000 387.650000 ;
      RECT 466.500000 386.350000 499.500000 387.650000 ;
      RECT 457.500000 386.350000 458.500000 387.650000 ;
      RECT 416.500000 386.350000 449.500000 387.650000 ;
      RECT 407.500000 386.350000 408.500000 387.650000 ;
      RECT 366.500000 386.350000 399.500000 387.650000 ;
      RECT 357.500000 386.350000 358.500000 387.650000 ;
      RECT 316.500000 386.350000 349.500000 387.650000 ;
      RECT 307.500000 386.350000 308.500000 387.650000 ;
      RECT 266.500000 386.350000 299.500000 387.650000 ;
      RECT 257.500000 386.350000 258.500000 387.650000 ;
      RECT 216.500000 386.350000 249.500000 387.650000 ;
      RECT 207.500000 386.350000 208.500000 387.650000 ;
      RECT 166.500000 386.350000 199.500000 387.650000 ;
      RECT 157.500000 386.350000 158.500000 387.650000 ;
      RECT 116.500000 386.350000 149.500000 387.650000 ;
      RECT 107.500000 386.350000 108.500000 387.650000 ;
      RECT 66.500000 386.350000 99.500000 387.650000 ;
      RECT 57.500000 386.350000 58.500000 387.650000 ;
      RECT 29.500000 386.350000 49.500000 387.650000 ;
      RECT 15.500000 386.350000 16.500000 387.650000 ;
      RECT 1157.500000 385.650000 1170.500000 386.350000 ;
      RECT 1107.500000 385.650000 1149.500000 386.350000 ;
      RECT 1057.500000 385.650000 1099.500000 386.350000 ;
      RECT 1007.500000 385.650000 1049.500000 386.350000 ;
      RECT 957.500000 385.650000 999.500000 386.350000 ;
      RECT 907.500000 385.650000 949.500000 386.350000 ;
      RECT 857.500000 385.650000 899.500000 386.350000 ;
      RECT 807.500000 385.650000 849.500000 386.350000 ;
      RECT 757.500000 385.650000 799.500000 386.350000 ;
      RECT 707.500000 385.650000 749.500000 386.350000 ;
      RECT 657.500000 385.650000 699.500000 386.350000 ;
      RECT 607.500000 385.650000 649.500000 386.350000 ;
      RECT 557.500000 385.650000 599.500000 386.350000 ;
      RECT 507.500000 385.650000 549.500000 386.350000 ;
      RECT 457.500000 385.650000 499.500000 386.350000 ;
      RECT 407.500000 385.650000 449.500000 386.350000 ;
      RECT 357.500000 385.650000 399.500000 386.350000 ;
      RECT 307.500000 385.650000 349.500000 386.350000 ;
      RECT 257.500000 385.650000 299.500000 386.350000 ;
      RECT 207.500000 385.650000 249.500000 386.350000 ;
      RECT 157.500000 385.650000 199.500000 386.350000 ;
      RECT 107.500000 385.650000 149.500000 386.350000 ;
      RECT 57.500000 385.650000 99.500000 386.350000 ;
      RECT 15.500000 385.650000 49.500000 386.350000 ;
      RECT 1183.500000 384.350000 1186.000000 387.650000 ;
      RECT 1169.500000 384.350000 1170.500000 385.650000 ;
      RECT 1116.500000 384.350000 1149.500000 385.650000 ;
      RECT 1107.500000 384.350000 1108.500000 385.650000 ;
      RECT 1066.500000 384.350000 1099.500000 385.650000 ;
      RECT 1057.500000 384.350000 1058.500000 385.650000 ;
      RECT 1016.500000 384.350000 1049.500000 385.650000 ;
      RECT 1007.500000 384.350000 1008.500000 385.650000 ;
      RECT 966.500000 384.350000 999.500000 385.650000 ;
      RECT 957.500000 384.350000 958.500000 385.650000 ;
      RECT 916.500000 384.350000 949.500000 385.650000 ;
      RECT 907.500000 384.350000 908.500000 385.650000 ;
      RECT 866.500000 384.350000 899.500000 385.650000 ;
      RECT 857.500000 384.350000 858.500000 385.650000 ;
      RECT 816.500000 384.350000 849.500000 385.650000 ;
      RECT 807.500000 384.350000 808.500000 385.650000 ;
      RECT 766.500000 384.350000 799.500000 385.650000 ;
      RECT 757.500000 384.350000 758.500000 385.650000 ;
      RECT 716.500000 384.350000 749.500000 385.650000 ;
      RECT 707.500000 384.350000 708.500000 385.650000 ;
      RECT 666.500000 384.350000 699.500000 385.650000 ;
      RECT 657.500000 384.350000 658.500000 385.650000 ;
      RECT 616.500000 384.350000 649.500000 385.650000 ;
      RECT 607.500000 384.350000 608.500000 385.650000 ;
      RECT 566.500000 384.350000 599.500000 385.650000 ;
      RECT 557.500000 384.350000 558.500000 385.650000 ;
      RECT 516.500000 384.350000 549.500000 385.650000 ;
      RECT 507.500000 384.350000 508.500000 385.650000 ;
      RECT 466.500000 384.350000 499.500000 385.650000 ;
      RECT 457.500000 384.350000 458.500000 385.650000 ;
      RECT 416.500000 384.350000 449.500000 385.650000 ;
      RECT 407.500000 384.350000 408.500000 385.650000 ;
      RECT 366.500000 384.350000 399.500000 385.650000 ;
      RECT 357.500000 384.350000 358.500000 385.650000 ;
      RECT 316.500000 384.350000 349.500000 385.650000 ;
      RECT 307.500000 384.350000 308.500000 385.650000 ;
      RECT 266.500000 384.350000 299.500000 385.650000 ;
      RECT 257.500000 384.350000 258.500000 385.650000 ;
      RECT 216.500000 384.350000 249.500000 385.650000 ;
      RECT 207.500000 384.350000 208.500000 385.650000 ;
      RECT 166.500000 384.350000 199.500000 385.650000 ;
      RECT 157.500000 384.350000 158.500000 385.650000 ;
      RECT 116.500000 384.350000 149.500000 385.650000 ;
      RECT 107.500000 384.350000 108.500000 385.650000 ;
      RECT 66.500000 384.350000 99.500000 385.650000 ;
      RECT 57.500000 384.350000 58.500000 385.650000 ;
      RECT 29.500000 384.350000 49.500000 385.650000 ;
      RECT 15.500000 384.350000 16.500000 385.650000 ;
      RECT 0.000000 384.350000 2.500000 387.650000 ;
      RECT 1169.500000 383.650000 1186.000000 384.350000 ;
      RECT 1116.500000 383.650000 1156.500000 384.350000 ;
      RECT 1066.500000 383.650000 1108.500000 384.350000 ;
      RECT 1016.500000 383.650000 1058.500000 384.350000 ;
      RECT 966.500000 383.650000 1008.500000 384.350000 ;
      RECT 916.500000 383.650000 958.500000 384.350000 ;
      RECT 866.500000 383.650000 908.500000 384.350000 ;
      RECT 816.500000 383.650000 858.500000 384.350000 ;
      RECT 766.500000 383.650000 808.500000 384.350000 ;
      RECT 716.500000 383.650000 758.500000 384.350000 ;
      RECT 666.500000 383.650000 708.500000 384.350000 ;
      RECT 616.500000 383.650000 658.500000 384.350000 ;
      RECT 566.500000 383.650000 608.500000 384.350000 ;
      RECT 516.500000 383.650000 558.500000 384.350000 ;
      RECT 466.500000 383.650000 508.500000 384.350000 ;
      RECT 416.500000 383.650000 458.500000 384.350000 ;
      RECT 366.500000 383.650000 408.500000 384.350000 ;
      RECT 316.500000 383.650000 358.500000 384.350000 ;
      RECT 266.500000 383.650000 308.500000 384.350000 ;
      RECT 216.500000 383.650000 258.500000 384.350000 ;
      RECT 166.500000 383.650000 208.500000 384.350000 ;
      RECT 116.500000 383.650000 158.500000 384.350000 ;
      RECT 66.500000 383.650000 108.500000 384.350000 ;
      RECT 29.500000 383.650000 58.500000 384.350000 ;
      RECT 0.000000 383.650000 16.500000 384.350000 ;
      RECT 1169.500000 382.350000 1170.500000 383.650000 ;
      RECT 1116.500000 382.350000 1149.500000 383.650000 ;
      RECT 1107.500000 382.350000 1108.500000 383.650000 ;
      RECT 1066.500000 382.350000 1099.500000 383.650000 ;
      RECT 1057.500000 382.350000 1058.500000 383.650000 ;
      RECT 1016.500000 382.350000 1049.500000 383.650000 ;
      RECT 1007.500000 382.350000 1008.500000 383.650000 ;
      RECT 966.500000 382.350000 999.500000 383.650000 ;
      RECT 957.500000 382.350000 958.500000 383.650000 ;
      RECT 916.500000 382.350000 949.500000 383.650000 ;
      RECT 907.500000 382.350000 908.500000 383.650000 ;
      RECT 866.500000 382.350000 899.500000 383.650000 ;
      RECT 857.500000 382.350000 858.500000 383.650000 ;
      RECT 816.500000 382.350000 849.500000 383.650000 ;
      RECT 807.500000 382.350000 808.500000 383.650000 ;
      RECT 766.500000 382.350000 799.500000 383.650000 ;
      RECT 757.500000 382.350000 758.500000 383.650000 ;
      RECT 716.500000 382.350000 749.500000 383.650000 ;
      RECT 707.500000 382.350000 708.500000 383.650000 ;
      RECT 666.500000 382.350000 699.500000 383.650000 ;
      RECT 657.500000 382.350000 658.500000 383.650000 ;
      RECT 616.500000 382.350000 649.500000 383.650000 ;
      RECT 607.500000 382.350000 608.500000 383.650000 ;
      RECT 566.500000 382.350000 599.500000 383.650000 ;
      RECT 557.500000 382.350000 558.500000 383.650000 ;
      RECT 516.500000 382.350000 549.500000 383.650000 ;
      RECT 507.500000 382.350000 508.500000 383.650000 ;
      RECT 466.500000 382.350000 499.500000 383.650000 ;
      RECT 457.500000 382.350000 458.500000 383.650000 ;
      RECT 416.500000 382.350000 449.500000 383.650000 ;
      RECT 407.500000 382.350000 408.500000 383.650000 ;
      RECT 366.500000 382.350000 399.500000 383.650000 ;
      RECT 357.500000 382.350000 358.500000 383.650000 ;
      RECT 316.500000 382.350000 349.500000 383.650000 ;
      RECT 307.500000 382.350000 308.500000 383.650000 ;
      RECT 266.500000 382.350000 299.500000 383.650000 ;
      RECT 257.500000 382.350000 258.500000 383.650000 ;
      RECT 216.500000 382.350000 249.500000 383.650000 ;
      RECT 207.500000 382.350000 208.500000 383.650000 ;
      RECT 166.500000 382.350000 199.500000 383.650000 ;
      RECT 157.500000 382.350000 158.500000 383.650000 ;
      RECT 116.500000 382.350000 149.500000 383.650000 ;
      RECT 107.500000 382.350000 108.500000 383.650000 ;
      RECT 66.500000 382.350000 99.500000 383.650000 ;
      RECT 57.500000 382.350000 58.500000 383.650000 ;
      RECT 29.500000 382.350000 49.500000 383.650000 ;
      RECT 15.500000 382.350000 16.500000 383.650000 ;
      RECT 1157.500000 381.650000 1170.500000 382.350000 ;
      RECT 1107.500000 381.650000 1149.500000 382.350000 ;
      RECT 1057.500000 381.650000 1099.500000 382.350000 ;
      RECT 1007.500000 381.650000 1049.500000 382.350000 ;
      RECT 957.500000 381.650000 999.500000 382.350000 ;
      RECT 907.500000 381.650000 949.500000 382.350000 ;
      RECT 857.500000 381.650000 899.500000 382.350000 ;
      RECT 807.500000 381.650000 849.500000 382.350000 ;
      RECT 757.500000 381.650000 799.500000 382.350000 ;
      RECT 707.500000 381.650000 749.500000 382.350000 ;
      RECT 657.500000 381.650000 699.500000 382.350000 ;
      RECT 607.500000 381.650000 649.500000 382.350000 ;
      RECT 557.500000 381.650000 599.500000 382.350000 ;
      RECT 507.500000 381.650000 549.500000 382.350000 ;
      RECT 457.500000 381.650000 499.500000 382.350000 ;
      RECT 407.500000 381.650000 449.500000 382.350000 ;
      RECT 357.500000 381.650000 399.500000 382.350000 ;
      RECT 307.500000 381.650000 349.500000 382.350000 ;
      RECT 257.500000 381.650000 299.500000 382.350000 ;
      RECT 207.500000 381.650000 249.500000 382.350000 ;
      RECT 157.500000 381.650000 199.500000 382.350000 ;
      RECT 107.500000 381.650000 149.500000 382.350000 ;
      RECT 57.500000 381.650000 99.500000 382.350000 ;
      RECT 15.500000 381.650000 49.500000 382.350000 ;
      RECT 1183.500000 380.350000 1186.000000 383.650000 ;
      RECT 1169.500000 380.350000 1170.500000 381.650000 ;
      RECT 1116.500000 380.350000 1149.500000 381.650000 ;
      RECT 1107.500000 380.350000 1108.500000 381.650000 ;
      RECT 1066.500000 380.350000 1099.500000 381.650000 ;
      RECT 1057.500000 380.350000 1058.500000 381.650000 ;
      RECT 1016.500000 380.350000 1049.500000 381.650000 ;
      RECT 1007.500000 380.350000 1008.500000 381.650000 ;
      RECT 966.500000 380.350000 999.500000 381.650000 ;
      RECT 957.500000 380.350000 958.500000 381.650000 ;
      RECT 916.500000 380.350000 949.500000 381.650000 ;
      RECT 907.500000 380.350000 908.500000 381.650000 ;
      RECT 866.500000 380.350000 899.500000 381.650000 ;
      RECT 857.500000 380.350000 858.500000 381.650000 ;
      RECT 816.500000 380.350000 849.500000 381.650000 ;
      RECT 807.500000 380.350000 808.500000 381.650000 ;
      RECT 766.500000 380.350000 799.500000 381.650000 ;
      RECT 757.500000 380.350000 758.500000 381.650000 ;
      RECT 716.500000 380.350000 749.500000 381.650000 ;
      RECT 707.500000 380.350000 708.500000 381.650000 ;
      RECT 666.500000 380.350000 699.500000 381.650000 ;
      RECT 657.500000 380.350000 658.500000 381.650000 ;
      RECT 616.500000 380.350000 649.500000 381.650000 ;
      RECT 607.500000 380.350000 608.500000 381.650000 ;
      RECT 566.500000 380.350000 599.500000 381.650000 ;
      RECT 557.500000 380.350000 558.500000 381.650000 ;
      RECT 516.500000 380.350000 549.500000 381.650000 ;
      RECT 507.500000 380.350000 508.500000 381.650000 ;
      RECT 466.500000 380.350000 499.500000 381.650000 ;
      RECT 457.500000 380.350000 458.500000 381.650000 ;
      RECT 416.500000 380.350000 449.500000 381.650000 ;
      RECT 407.500000 380.350000 408.500000 381.650000 ;
      RECT 366.500000 380.350000 399.500000 381.650000 ;
      RECT 357.500000 380.350000 358.500000 381.650000 ;
      RECT 316.500000 380.350000 349.500000 381.650000 ;
      RECT 307.500000 380.350000 308.500000 381.650000 ;
      RECT 266.500000 380.350000 299.500000 381.650000 ;
      RECT 257.500000 380.350000 258.500000 381.650000 ;
      RECT 216.500000 380.350000 249.500000 381.650000 ;
      RECT 207.500000 380.350000 208.500000 381.650000 ;
      RECT 166.500000 380.350000 199.500000 381.650000 ;
      RECT 157.500000 380.350000 158.500000 381.650000 ;
      RECT 116.500000 380.350000 149.500000 381.650000 ;
      RECT 107.500000 380.350000 108.500000 381.650000 ;
      RECT 66.500000 380.350000 99.500000 381.650000 ;
      RECT 57.500000 380.350000 58.500000 381.650000 ;
      RECT 29.500000 380.350000 49.500000 381.650000 ;
      RECT 15.500000 380.350000 16.500000 381.650000 ;
      RECT 0.000000 380.350000 2.500000 383.650000 ;
      RECT 1169.500000 379.650000 1186.000000 380.350000 ;
      RECT 1116.500000 379.650000 1156.500000 380.350000 ;
      RECT 1066.500000 379.650000 1108.500000 380.350000 ;
      RECT 1016.500000 379.650000 1058.500000 380.350000 ;
      RECT 966.500000 379.650000 1008.500000 380.350000 ;
      RECT 916.500000 379.650000 958.500000 380.350000 ;
      RECT 866.500000 379.650000 908.500000 380.350000 ;
      RECT 816.500000 379.650000 858.500000 380.350000 ;
      RECT 766.500000 379.650000 808.500000 380.350000 ;
      RECT 716.500000 379.650000 758.500000 380.350000 ;
      RECT 666.500000 379.650000 708.500000 380.350000 ;
      RECT 616.500000 379.650000 658.500000 380.350000 ;
      RECT 566.500000 379.650000 608.500000 380.350000 ;
      RECT 516.500000 379.650000 558.500000 380.350000 ;
      RECT 466.500000 379.650000 508.500000 380.350000 ;
      RECT 416.500000 379.650000 458.500000 380.350000 ;
      RECT 366.500000 379.650000 408.500000 380.350000 ;
      RECT 316.500000 379.650000 358.500000 380.350000 ;
      RECT 266.500000 379.650000 308.500000 380.350000 ;
      RECT 216.500000 379.650000 258.500000 380.350000 ;
      RECT 166.500000 379.650000 208.500000 380.350000 ;
      RECT 116.500000 379.650000 158.500000 380.350000 ;
      RECT 66.500000 379.650000 108.500000 380.350000 ;
      RECT 29.500000 379.650000 58.500000 380.350000 ;
      RECT 0.000000 379.650000 16.500000 380.350000 ;
      RECT 1169.500000 378.350000 1170.500000 379.650000 ;
      RECT 1116.500000 378.350000 1149.500000 379.650000 ;
      RECT 1107.500000 378.350000 1108.500000 379.650000 ;
      RECT 1066.500000 378.350000 1099.500000 379.650000 ;
      RECT 1057.500000 378.350000 1058.500000 379.650000 ;
      RECT 1016.500000 378.350000 1049.500000 379.650000 ;
      RECT 1007.500000 378.350000 1008.500000 379.650000 ;
      RECT 966.500000 378.350000 999.500000 379.650000 ;
      RECT 957.500000 378.350000 958.500000 379.650000 ;
      RECT 916.500000 378.350000 949.500000 379.650000 ;
      RECT 907.500000 378.350000 908.500000 379.650000 ;
      RECT 866.500000 378.350000 899.500000 379.650000 ;
      RECT 857.500000 378.350000 858.500000 379.650000 ;
      RECT 816.500000 378.350000 849.500000 379.650000 ;
      RECT 807.500000 378.350000 808.500000 379.650000 ;
      RECT 766.500000 378.350000 799.500000 379.650000 ;
      RECT 757.500000 378.350000 758.500000 379.650000 ;
      RECT 716.500000 378.350000 749.500000 379.650000 ;
      RECT 707.500000 378.350000 708.500000 379.650000 ;
      RECT 666.500000 378.350000 699.500000 379.650000 ;
      RECT 657.500000 378.350000 658.500000 379.650000 ;
      RECT 616.500000 378.350000 649.500000 379.650000 ;
      RECT 607.500000 378.350000 608.500000 379.650000 ;
      RECT 566.500000 378.350000 599.500000 379.650000 ;
      RECT 557.500000 378.350000 558.500000 379.650000 ;
      RECT 516.500000 378.350000 549.500000 379.650000 ;
      RECT 507.500000 378.350000 508.500000 379.650000 ;
      RECT 466.500000 378.350000 499.500000 379.650000 ;
      RECT 457.500000 378.350000 458.500000 379.650000 ;
      RECT 416.500000 378.350000 449.500000 379.650000 ;
      RECT 407.500000 378.350000 408.500000 379.650000 ;
      RECT 366.500000 378.350000 399.500000 379.650000 ;
      RECT 357.500000 378.350000 358.500000 379.650000 ;
      RECT 316.500000 378.350000 349.500000 379.650000 ;
      RECT 307.500000 378.350000 308.500000 379.650000 ;
      RECT 266.500000 378.350000 299.500000 379.650000 ;
      RECT 257.500000 378.350000 258.500000 379.650000 ;
      RECT 216.500000 378.350000 249.500000 379.650000 ;
      RECT 207.500000 378.350000 208.500000 379.650000 ;
      RECT 166.500000 378.350000 199.500000 379.650000 ;
      RECT 157.500000 378.350000 158.500000 379.650000 ;
      RECT 116.500000 378.350000 149.500000 379.650000 ;
      RECT 107.500000 378.350000 108.500000 379.650000 ;
      RECT 66.500000 378.350000 99.500000 379.650000 ;
      RECT 57.500000 378.350000 58.500000 379.650000 ;
      RECT 29.500000 378.350000 49.500000 379.650000 ;
      RECT 15.500000 378.350000 16.500000 379.650000 ;
      RECT 1157.500000 377.650000 1170.500000 378.350000 ;
      RECT 1107.500000 377.650000 1149.500000 378.350000 ;
      RECT 1057.500000 377.650000 1099.500000 378.350000 ;
      RECT 1007.500000 377.650000 1049.500000 378.350000 ;
      RECT 957.500000 377.650000 999.500000 378.350000 ;
      RECT 907.500000 377.650000 949.500000 378.350000 ;
      RECT 857.500000 377.650000 899.500000 378.350000 ;
      RECT 807.500000 377.650000 849.500000 378.350000 ;
      RECT 757.500000 377.650000 799.500000 378.350000 ;
      RECT 707.500000 377.650000 749.500000 378.350000 ;
      RECT 657.500000 377.650000 699.500000 378.350000 ;
      RECT 607.500000 377.650000 649.500000 378.350000 ;
      RECT 557.500000 377.650000 599.500000 378.350000 ;
      RECT 507.500000 377.650000 549.500000 378.350000 ;
      RECT 457.500000 377.650000 499.500000 378.350000 ;
      RECT 407.500000 377.650000 449.500000 378.350000 ;
      RECT 357.500000 377.650000 399.500000 378.350000 ;
      RECT 307.500000 377.650000 349.500000 378.350000 ;
      RECT 257.500000 377.650000 299.500000 378.350000 ;
      RECT 207.500000 377.650000 249.500000 378.350000 ;
      RECT 157.500000 377.650000 199.500000 378.350000 ;
      RECT 107.500000 377.650000 149.500000 378.350000 ;
      RECT 57.500000 377.650000 99.500000 378.350000 ;
      RECT 15.500000 377.650000 49.500000 378.350000 ;
      RECT 1183.500000 376.350000 1186.000000 379.650000 ;
      RECT 1169.500000 376.350000 1170.500000 377.650000 ;
      RECT 1116.500000 376.350000 1149.500000 377.650000 ;
      RECT 1107.500000 376.350000 1108.500000 377.650000 ;
      RECT 1066.500000 376.350000 1099.500000 377.650000 ;
      RECT 1057.500000 376.350000 1058.500000 377.650000 ;
      RECT 1016.500000 376.350000 1049.500000 377.650000 ;
      RECT 1007.500000 376.350000 1008.500000 377.650000 ;
      RECT 966.500000 376.350000 999.500000 377.650000 ;
      RECT 957.500000 376.350000 958.500000 377.650000 ;
      RECT 916.500000 376.350000 949.500000 377.650000 ;
      RECT 907.500000 376.350000 908.500000 377.650000 ;
      RECT 866.500000 376.350000 899.500000 377.650000 ;
      RECT 857.500000 376.350000 858.500000 377.650000 ;
      RECT 816.500000 376.350000 849.500000 377.650000 ;
      RECT 807.500000 376.350000 808.500000 377.650000 ;
      RECT 766.500000 376.350000 799.500000 377.650000 ;
      RECT 757.500000 376.350000 758.500000 377.650000 ;
      RECT 716.500000 376.350000 749.500000 377.650000 ;
      RECT 707.500000 376.350000 708.500000 377.650000 ;
      RECT 666.500000 376.350000 699.500000 377.650000 ;
      RECT 657.500000 376.350000 658.500000 377.650000 ;
      RECT 616.500000 376.350000 649.500000 377.650000 ;
      RECT 607.500000 376.350000 608.500000 377.650000 ;
      RECT 566.500000 376.350000 599.500000 377.650000 ;
      RECT 557.500000 376.350000 558.500000 377.650000 ;
      RECT 516.500000 376.350000 549.500000 377.650000 ;
      RECT 507.500000 376.350000 508.500000 377.650000 ;
      RECT 466.500000 376.350000 499.500000 377.650000 ;
      RECT 457.500000 376.350000 458.500000 377.650000 ;
      RECT 416.500000 376.350000 449.500000 377.650000 ;
      RECT 407.500000 376.350000 408.500000 377.650000 ;
      RECT 366.500000 376.350000 399.500000 377.650000 ;
      RECT 357.500000 376.350000 358.500000 377.650000 ;
      RECT 316.500000 376.350000 349.500000 377.650000 ;
      RECT 307.500000 376.350000 308.500000 377.650000 ;
      RECT 266.500000 376.350000 299.500000 377.650000 ;
      RECT 257.500000 376.350000 258.500000 377.650000 ;
      RECT 216.500000 376.350000 249.500000 377.650000 ;
      RECT 207.500000 376.350000 208.500000 377.650000 ;
      RECT 166.500000 376.350000 199.500000 377.650000 ;
      RECT 157.500000 376.350000 158.500000 377.650000 ;
      RECT 116.500000 376.350000 149.500000 377.650000 ;
      RECT 107.500000 376.350000 108.500000 377.650000 ;
      RECT 66.500000 376.350000 99.500000 377.650000 ;
      RECT 57.500000 376.350000 58.500000 377.650000 ;
      RECT 29.500000 376.350000 49.500000 377.650000 ;
      RECT 15.500000 376.350000 16.500000 377.650000 ;
      RECT 0.000000 376.350000 2.500000 379.650000 ;
      RECT 1169.500000 375.650000 1186.000000 376.350000 ;
      RECT 1116.500000 375.650000 1156.500000 376.350000 ;
      RECT 1066.500000 375.650000 1108.500000 376.350000 ;
      RECT 1016.500000 375.650000 1058.500000 376.350000 ;
      RECT 966.500000 375.650000 1008.500000 376.350000 ;
      RECT 916.500000 375.650000 958.500000 376.350000 ;
      RECT 866.500000 375.650000 908.500000 376.350000 ;
      RECT 816.500000 375.650000 858.500000 376.350000 ;
      RECT 766.500000 375.650000 808.500000 376.350000 ;
      RECT 716.500000 375.650000 758.500000 376.350000 ;
      RECT 666.500000 375.650000 708.500000 376.350000 ;
      RECT 616.500000 375.650000 658.500000 376.350000 ;
      RECT 566.500000 375.650000 608.500000 376.350000 ;
      RECT 516.500000 375.650000 558.500000 376.350000 ;
      RECT 466.500000 375.650000 508.500000 376.350000 ;
      RECT 416.500000 375.650000 458.500000 376.350000 ;
      RECT 366.500000 375.650000 408.500000 376.350000 ;
      RECT 316.500000 375.650000 358.500000 376.350000 ;
      RECT 266.500000 375.650000 308.500000 376.350000 ;
      RECT 216.500000 375.650000 258.500000 376.350000 ;
      RECT 166.500000 375.650000 208.500000 376.350000 ;
      RECT 116.500000 375.650000 158.500000 376.350000 ;
      RECT 66.500000 375.650000 108.500000 376.350000 ;
      RECT 29.500000 375.650000 58.500000 376.350000 ;
      RECT 0.000000 375.650000 16.500000 376.350000 ;
      RECT 1169.500000 374.350000 1170.500000 375.650000 ;
      RECT 1116.500000 374.350000 1149.500000 375.650000 ;
      RECT 1107.500000 374.350000 1108.500000 375.650000 ;
      RECT 1066.500000 374.350000 1099.500000 375.650000 ;
      RECT 1057.500000 374.350000 1058.500000 375.650000 ;
      RECT 1016.500000 374.350000 1049.500000 375.650000 ;
      RECT 1007.500000 374.350000 1008.500000 375.650000 ;
      RECT 966.500000 374.350000 999.500000 375.650000 ;
      RECT 957.500000 374.350000 958.500000 375.650000 ;
      RECT 916.500000 374.350000 949.500000 375.650000 ;
      RECT 907.500000 374.350000 908.500000 375.650000 ;
      RECT 866.500000 374.350000 899.500000 375.650000 ;
      RECT 857.500000 374.350000 858.500000 375.650000 ;
      RECT 816.500000 374.350000 849.500000 375.650000 ;
      RECT 807.500000 374.350000 808.500000 375.650000 ;
      RECT 766.500000 374.350000 799.500000 375.650000 ;
      RECT 757.500000 374.350000 758.500000 375.650000 ;
      RECT 716.500000 374.350000 749.500000 375.650000 ;
      RECT 707.500000 374.350000 708.500000 375.650000 ;
      RECT 666.500000 374.350000 699.500000 375.650000 ;
      RECT 657.500000 374.350000 658.500000 375.650000 ;
      RECT 616.500000 374.350000 649.500000 375.650000 ;
      RECT 607.500000 374.350000 608.500000 375.650000 ;
      RECT 566.500000 374.350000 599.500000 375.650000 ;
      RECT 557.500000 374.350000 558.500000 375.650000 ;
      RECT 516.500000 374.350000 549.500000 375.650000 ;
      RECT 507.500000 374.350000 508.500000 375.650000 ;
      RECT 466.500000 374.350000 499.500000 375.650000 ;
      RECT 457.500000 374.350000 458.500000 375.650000 ;
      RECT 416.500000 374.350000 449.500000 375.650000 ;
      RECT 407.500000 374.350000 408.500000 375.650000 ;
      RECT 366.500000 374.350000 399.500000 375.650000 ;
      RECT 357.500000 374.350000 358.500000 375.650000 ;
      RECT 316.500000 374.350000 349.500000 375.650000 ;
      RECT 307.500000 374.350000 308.500000 375.650000 ;
      RECT 266.500000 374.350000 299.500000 375.650000 ;
      RECT 257.500000 374.350000 258.500000 375.650000 ;
      RECT 216.500000 374.350000 249.500000 375.650000 ;
      RECT 207.500000 374.350000 208.500000 375.650000 ;
      RECT 166.500000 374.350000 199.500000 375.650000 ;
      RECT 157.500000 374.350000 158.500000 375.650000 ;
      RECT 116.500000 374.350000 149.500000 375.650000 ;
      RECT 107.500000 374.350000 108.500000 375.650000 ;
      RECT 66.500000 374.350000 99.500000 375.650000 ;
      RECT 57.500000 374.350000 58.500000 375.650000 ;
      RECT 29.500000 374.350000 49.500000 375.650000 ;
      RECT 15.500000 374.350000 16.500000 375.650000 ;
      RECT 1157.500000 373.650000 1170.500000 374.350000 ;
      RECT 1107.500000 373.650000 1149.500000 374.350000 ;
      RECT 1057.500000 373.650000 1099.500000 374.350000 ;
      RECT 1007.500000 373.650000 1049.500000 374.350000 ;
      RECT 957.500000 373.650000 999.500000 374.350000 ;
      RECT 907.500000 373.650000 949.500000 374.350000 ;
      RECT 857.500000 373.650000 899.500000 374.350000 ;
      RECT 807.500000 373.650000 849.500000 374.350000 ;
      RECT 757.500000 373.650000 799.500000 374.350000 ;
      RECT 707.500000 373.650000 749.500000 374.350000 ;
      RECT 657.500000 373.650000 699.500000 374.350000 ;
      RECT 607.500000 373.650000 649.500000 374.350000 ;
      RECT 557.500000 373.650000 599.500000 374.350000 ;
      RECT 507.500000 373.650000 549.500000 374.350000 ;
      RECT 457.500000 373.650000 499.500000 374.350000 ;
      RECT 407.500000 373.650000 449.500000 374.350000 ;
      RECT 357.500000 373.650000 399.500000 374.350000 ;
      RECT 307.500000 373.650000 349.500000 374.350000 ;
      RECT 257.500000 373.650000 299.500000 374.350000 ;
      RECT 207.500000 373.650000 249.500000 374.350000 ;
      RECT 157.500000 373.650000 199.500000 374.350000 ;
      RECT 107.500000 373.650000 149.500000 374.350000 ;
      RECT 57.500000 373.650000 99.500000 374.350000 ;
      RECT 15.500000 373.650000 49.500000 374.350000 ;
      RECT 1183.500000 372.350000 1186.000000 375.650000 ;
      RECT 1169.500000 372.350000 1170.500000 373.650000 ;
      RECT 1116.500000 372.350000 1149.500000 373.650000 ;
      RECT 1107.500000 372.350000 1108.500000 373.650000 ;
      RECT 1066.500000 372.350000 1099.500000 373.650000 ;
      RECT 1057.500000 372.350000 1058.500000 373.650000 ;
      RECT 1016.500000 372.350000 1049.500000 373.650000 ;
      RECT 1007.500000 372.350000 1008.500000 373.650000 ;
      RECT 966.500000 372.350000 999.500000 373.650000 ;
      RECT 957.500000 372.350000 958.500000 373.650000 ;
      RECT 916.500000 372.350000 949.500000 373.650000 ;
      RECT 907.500000 372.350000 908.500000 373.650000 ;
      RECT 866.500000 372.350000 899.500000 373.650000 ;
      RECT 857.500000 372.350000 858.500000 373.650000 ;
      RECT 816.500000 372.350000 849.500000 373.650000 ;
      RECT 807.500000 372.350000 808.500000 373.650000 ;
      RECT 766.500000 372.350000 799.500000 373.650000 ;
      RECT 757.500000 372.350000 758.500000 373.650000 ;
      RECT 716.500000 372.350000 749.500000 373.650000 ;
      RECT 707.500000 372.350000 708.500000 373.650000 ;
      RECT 666.500000 372.350000 699.500000 373.650000 ;
      RECT 657.500000 372.350000 658.500000 373.650000 ;
      RECT 616.500000 372.350000 649.500000 373.650000 ;
      RECT 607.500000 372.350000 608.500000 373.650000 ;
      RECT 566.500000 372.350000 599.500000 373.650000 ;
      RECT 557.500000 372.350000 558.500000 373.650000 ;
      RECT 516.500000 372.350000 549.500000 373.650000 ;
      RECT 507.500000 372.350000 508.500000 373.650000 ;
      RECT 466.500000 372.350000 499.500000 373.650000 ;
      RECT 457.500000 372.350000 458.500000 373.650000 ;
      RECT 416.500000 372.350000 449.500000 373.650000 ;
      RECT 407.500000 372.350000 408.500000 373.650000 ;
      RECT 366.500000 372.350000 399.500000 373.650000 ;
      RECT 357.500000 372.350000 358.500000 373.650000 ;
      RECT 316.500000 372.350000 349.500000 373.650000 ;
      RECT 307.500000 372.350000 308.500000 373.650000 ;
      RECT 266.500000 372.350000 299.500000 373.650000 ;
      RECT 257.500000 372.350000 258.500000 373.650000 ;
      RECT 216.500000 372.350000 249.500000 373.650000 ;
      RECT 207.500000 372.350000 208.500000 373.650000 ;
      RECT 166.500000 372.350000 199.500000 373.650000 ;
      RECT 157.500000 372.350000 158.500000 373.650000 ;
      RECT 116.500000 372.350000 149.500000 373.650000 ;
      RECT 107.500000 372.350000 108.500000 373.650000 ;
      RECT 66.500000 372.350000 99.500000 373.650000 ;
      RECT 57.500000 372.350000 58.500000 373.650000 ;
      RECT 29.500000 372.350000 49.500000 373.650000 ;
      RECT 15.500000 372.350000 16.500000 373.650000 ;
      RECT 0.000000 372.350000 2.500000 375.650000 ;
      RECT 1169.500000 371.650000 1186.000000 372.350000 ;
      RECT 1116.500000 371.650000 1156.500000 372.350000 ;
      RECT 1066.500000 371.650000 1108.500000 372.350000 ;
      RECT 1016.500000 371.650000 1058.500000 372.350000 ;
      RECT 966.500000 371.650000 1008.500000 372.350000 ;
      RECT 916.500000 371.650000 958.500000 372.350000 ;
      RECT 866.500000 371.650000 908.500000 372.350000 ;
      RECT 816.500000 371.650000 858.500000 372.350000 ;
      RECT 766.500000 371.650000 808.500000 372.350000 ;
      RECT 716.500000 371.650000 758.500000 372.350000 ;
      RECT 666.500000 371.650000 708.500000 372.350000 ;
      RECT 616.500000 371.650000 658.500000 372.350000 ;
      RECT 566.500000 371.650000 608.500000 372.350000 ;
      RECT 516.500000 371.650000 558.500000 372.350000 ;
      RECT 466.500000 371.650000 508.500000 372.350000 ;
      RECT 416.500000 371.650000 458.500000 372.350000 ;
      RECT 366.500000 371.650000 408.500000 372.350000 ;
      RECT 316.500000 371.650000 358.500000 372.350000 ;
      RECT 266.500000 371.650000 308.500000 372.350000 ;
      RECT 216.500000 371.650000 258.500000 372.350000 ;
      RECT 166.500000 371.650000 208.500000 372.350000 ;
      RECT 116.500000 371.650000 158.500000 372.350000 ;
      RECT 66.500000 371.650000 108.500000 372.350000 ;
      RECT 29.500000 371.650000 58.500000 372.350000 ;
      RECT 0.000000 371.650000 16.500000 372.350000 ;
      RECT 1169.500000 370.350000 1170.500000 371.650000 ;
      RECT 1116.500000 370.350000 1149.500000 371.650000 ;
      RECT 1107.500000 370.350000 1108.500000 371.650000 ;
      RECT 1066.500000 370.350000 1099.500000 371.650000 ;
      RECT 1057.500000 370.350000 1058.500000 371.650000 ;
      RECT 1016.500000 370.350000 1049.500000 371.650000 ;
      RECT 1007.500000 370.350000 1008.500000 371.650000 ;
      RECT 966.500000 370.350000 999.500000 371.650000 ;
      RECT 957.500000 370.350000 958.500000 371.650000 ;
      RECT 916.500000 370.350000 949.500000 371.650000 ;
      RECT 907.500000 370.350000 908.500000 371.650000 ;
      RECT 866.500000 370.350000 899.500000 371.650000 ;
      RECT 857.500000 370.350000 858.500000 371.650000 ;
      RECT 816.500000 370.350000 849.500000 371.650000 ;
      RECT 807.500000 370.350000 808.500000 371.650000 ;
      RECT 766.500000 370.350000 799.500000 371.650000 ;
      RECT 757.500000 370.350000 758.500000 371.650000 ;
      RECT 716.500000 370.350000 749.500000 371.650000 ;
      RECT 707.500000 370.350000 708.500000 371.650000 ;
      RECT 666.500000 370.350000 699.500000 371.650000 ;
      RECT 657.500000 370.350000 658.500000 371.650000 ;
      RECT 616.500000 370.350000 649.500000 371.650000 ;
      RECT 607.500000 370.350000 608.500000 371.650000 ;
      RECT 566.500000 370.350000 599.500000 371.650000 ;
      RECT 557.500000 370.350000 558.500000 371.650000 ;
      RECT 516.500000 370.350000 549.500000 371.650000 ;
      RECT 507.500000 370.350000 508.500000 371.650000 ;
      RECT 466.500000 370.350000 499.500000 371.650000 ;
      RECT 457.500000 370.350000 458.500000 371.650000 ;
      RECT 416.500000 370.350000 449.500000 371.650000 ;
      RECT 407.500000 370.350000 408.500000 371.650000 ;
      RECT 366.500000 370.350000 399.500000 371.650000 ;
      RECT 357.500000 370.350000 358.500000 371.650000 ;
      RECT 316.500000 370.350000 349.500000 371.650000 ;
      RECT 307.500000 370.350000 308.500000 371.650000 ;
      RECT 266.500000 370.350000 299.500000 371.650000 ;
      RECT 257.500000 370.350000 258.500000 371.650000 ;
      RECT 216.500000 370.350000 249.500000 371.650000 ;
      RECT 207.500000 370.350000 208.500000 371.650000 ;
      RECT 166.500000 370.350000 199.500000 371.650000 ;
      RECT 157.500000 370.350000 158.500000 371.650000 ;
      RECT 116.500000 370.350000 149.500000 371.650000 ;
      RECT 107.500000 370.350000 108.500000 371.650000 ;
      RECT 66.500000 370.350000 99.500000 371.650000 ;
      RECT 57.500000 370.350000 58.500000 371.650000 ;
      RECT 29.500000 370.350000 49.500000 371.650000 ;
      RECT 15.500000 370.350000 16.500000 371.650000 ;
      RECT 1157.500000 369.650000 1170.500000 370.350000 ;
      RECT 1107.500000 369.650000 1149.500000 370.350000 ;
      RECT 1057.500000 369.650000 1099.500000 370.350000 ;
      RECT 1007.500000 369.650000 1049.500000 370.350000 ;
      RECT 957.500000 369.650000 999.500000 370.350000 ;
      RECT 907.500000 369.650000 949.500000 370.350000 ;
      RECT 857.500000 369.650000 899.500000 370.350000 ;
      RECT 807.500000 369.650000 849.500000 370.350000 ;
      RECT 757.500000 369.650000 799.500000 370.350000 ;
      RECT 707.500000 369.650000 749.500000 370.350000 ;
      RECT 657.500000 369.650000 699.500000 370.350000 ;
      RECT 607.500000 369.650000 649.500000 370.350000 ;
      RECT 557.500000 369.650000 599.500000 370.350000 ;
      RECT 507.500000 369.650000 549.500000 370.350000 ;
      RECT 407.500000 369.650000 449.500000 370.350000 ;
      RECT 357.500000 369.650000 399.500000 370.350000 ;
      RECT 307.500000 369.650000 349.500000 370.350000 ;
      RECT 257.500000 369.650000 299.500000 370.350000 ;
      RECT 207.500000 369.650000 249.500000 370.350000 ;
      RECT 157.500000 369.650000 199.500000 370.350000 ;
      RECT 107.500000 369.650000 149.500000 370.350000 ;
      RECT 57.500000 369.650000 99.500000 370.350000 ;
      RECT 15.500000 369.650000 49.500000 370.350000 ;
      RECT 1183.500000 368.350000 1186.000000 371.650000 ;
      RECT 1169.500000 368.350000 1170.500000 369.650000 ;
      RECT 1116.500000 368.350000 1149.500000 369.650000 ;
      RECT 1107.500000 368.350000 1108.500000 369.650000 ;
      RECT 1066.500000 368.350000 1099.500000 369.650000 ;
      RECT 1057.500000 368.350000 1058.500000 369.650000 ;
      RECT 1016.500000 368.350000 1049.500000 369.650000 ;
      RECT 1007.500000 368.350000 1008.500000 369.650000 ;
      RECT 966.500000 368.350000 999.500000 369.650000 ;
      RECT 957.500000 368.350000 958.500000 369.650000 ;
      RECT 916.500000 368.350000 949.500000 369.650000 ;
      RECT 907.500000 368.350000 908.500000 369.650000 ;
      RECT 866.500000 368.350000 899.500000 369.650000 ;
      RECT 857.500000 368.350000 858.500000 369.650000 ;
      RECT 816.500000 368.350000 849.500000 369.650000 ;
      RECT 807.500000 368.350000 808.500000 369.650000 ;
      RECT 766.500000 368.350000 799.500000 369.650000 ;
      RECT 757.500000 368.350000 758.500000 369.650000 ;
      RECT 716.500000 368.350000 749.500000 369.650000 ;
      RECT 707.500000 368.350000 708.500000 369.650000 ;
      RECT 666.500000 368.350000 699.500000 369.650000 ;
      RECT 657.500000 368.350000 658.500000 369.650000 ;
      RECT 616.500000 368.350000 649.500000 369.650000 ;
      RECT 607.500000 368.350000 608.500000 369.650000 ;
      RECT 566.500000 368.350000 599.500000 369.650000 ;
      RECT 557.500000 368.350000 558.500000 369.650000 ;
      RECT 516.500000 368.350000 549.500000 369.650000 ;
      RECT 507.500000 368.350000 508.500000 369.650000 ;
      RECT 457.500000 368.350000 499.500000 370.350000 ;
      RECT 407.500000 368.350000 408.500000 369.650000 ;
      RECT 366.500000 368.350000 399.500000 369.650000 ;
      RECT 357.500000 368.350000 358.500000 369.650000 ;
      RECT 316.500000 368.350000 349.500000 369.650000 ;
      RECT 307.500000 368.350000 308.500000 369.650000 ;
      RECT 266.500000 368.350000 299.500000 369.650000 ;
      RECT 257.500000 368.350000 258.500000 369.650000 ;
      RECT 216.500000 368.350000 249.500000 369.650000 ;
      RECT 207.500000 368.350000 208.500000 369.650000 ;
      RECT 166.500000 368.350000 199.500000 369.650000 ;
      RECT 157.500000 368.350000 158.500000 369.650000 ;
      RECT 116.500000 368.350000 149.500000 369.650000 ;
      RECT 107.500000 368.350000 108.500000 369.650000 ;
      RECT 66.500000 368.350000 99.500000 369.650000 ;
      RECT 57.500000 368.350000 58.500000 369.650000 ;
      RECT 29.500000 368.350000 49.500000 369.650000 ;
      RECT 15.500000 368.350000 16.500000 369.650000 ;
      RECT 0.000000 368.350000 2.500000 371.650000 ;
      RECT 1169.500000 367.650000 1186.000000 368.350000 ;
      RECT 1116.500000 367.650000 1156.500000 368.350000 ;
      RECT 1066.500000 367.650000 1108.500000 368.350000 ;
      RECT 1016.500000 367.650000 1058.500000 368.350000 ;
      RECT 966.500000 367.650000 1008.500000 368.350000 ;
      RECT 916.500000 367.650000 958.500000 368.350000 ;
      RECT 866.500000 367.650000 908.500000 368.350000 ;
      RECT 816.500000 367.650000 858.500000 368.350000 ;
      RECT 766.500000 367.650000 808.500000 368.350000 ;
      RECT 716.500000 367.650000 758.500000 368.350000 ;
      RECT 666.500000 367.650000 708.500000 368.350000 ;
      RECT 616.500000 367.650000 658.500000 368.350000 ;
      RECT 566.500000 367.650000 608.500000 368.350000 ;
      RECT 516.500000 367.650000 558.500000 368.350000 ;
      RECT 457.500000 367.650000 508.500000 368.350000 ;
      RECT 366.500000 367.650000 408.500000 368.350000 ;
      RECT 316.500000 367.650000 358.500000 368.350000 ;
      RECT 266.500000 367.650000 308.500000 368.350000 ;
      RECT 216.500000 367.650000 258.500000 368.350000 ;
      RECT 166.500000 367.650000 208.500000 368.350000 ;
      RECT 116.500000 367.650000 158.500000 368.350000 ;
      RECT 66.500000 367.650000 108.500000 368.350000 ;
      RECT 29.500000 367.650000 58.500000 368.350000 ;
      RECT 0.000000 367.650000 16.500000 368.350000 ;
      RECT 1169.500000 366.350000 1170.500000 367.650000 ;
      RECT 1116.500000 366.350000 1149.500000 367.650000 ;
      RECT 1107.500000 366.350000 1108.500000 367.650000 ;
      RECT 1066.500000 366.350000 1099.500000 367.650000 ;
      RECT 1057.500000 366.350000 1058.500000 367.650000 ;
      RECT 1016.500000 366.350000 1049.500000 367.650000 ;
      RECT 1007.500000 366.350000 1008.500000 367.650000 ;
      RECT 966.500000 366.350000 999.500000 367.650000 ;
      RECT 957.500000 366.350000 958.500000 367.650000 ;
      RECT 916.500000 366.350000 949.500000 367.650000 ;
      RECT 907.500000 366.350000 908.500000 367.650000 ;
      RECT 866.500000 366.350000 899.500000 367.650000 ;
      RECT 857.500000 366.350000 858.500000 367.650000 ;
      RECT 816.500000 366.350000 849.500000 367.650000 ;
      RECT 807.500000 366.350000 808.500000 367.650000 ;
      RECT 766.500000 366.350000 799.500000 367.650000 ;
      RECT 757.500000 366.350000 758.500000 367.650000 ;
      RECT 716.500000 366.350000 749.500000 367.650000 ;
      RECT 707.500000 366.350000 708.500000 367.650000 ;
      RECT 666.500000 366.350000 699.500000 367.650000 ;
      RECT 657.500000 366.350000 658.500000 367.650000 ;
      RECT 616.500000 366.350000 649.500000 367.650000 ;
      RECT 607.500000 366.350000 608.500000 367.650000 ;
      RECT 566.500000 366.350000 599.500000 367.650000 ;
      RECT 557.500000 366.350000 558.500000 367.650000 ;
      RECT 516.500000 366.350000 549.500000 367.650000 ;
      RECT 507.500000 366.350000 508.500000 367.650000 ;
      RECT 416.500000 366.350000 449.500000 369.650000 ;
      RECT 407.500000 366.350000 408.500000 367.650000 ;
      RECT 366.500000 366.350000 399.500000 367.650000 ;
      RECT 357.500000 366.350000 358.500000 367.650000 ;
      RECT 316.500000 366.350000 349.500000 367.650000 ;
      RECT 307.500000 366.350000 308.500000 367.650000 ;
      RECT 266.500000 366.350000 299.500000 367.650000 ;
      RECT 257.500000 366.350000 258.500000 367.650000 ;
      RECT 216.500000 366.350000 249.500000 367.650000 ;
      RECT 207.500000 366.350000 208.500000 367.650000 ;
      RECT 166.500000 366.350000 199.500000 367.650000 ;
      RECT 157.500000 366.350000 158.500000 367.650000 ;
      RECT 116.500000 366.350000 149.500000 367.650000 ;
      RECT 107.500000 366.350000 108.500000 367.650000 ;
      RECT 66.500000 366.350000 99.500000 367.650000 ;
      RECT 57.500000 366.350000 58.500000 367.650000 ;
      RECT 29.500000 366.350000 49.500000 367.650000 ;
      RECT 15.500000 366.350000 16.500000 367.650000 ;
      RECT 1157.500000 365.650000 1170.500000 366.350000 ;
      RECT 1107.500000 365.650000 1149.500000 366.350000 ;
      RECT 1057.500000 365.650000 1099.500000 366.350000 ;
      RECT 1007.500000 365.650000 1049.500000 366.350000 ;
      RECT 957.500000 365.650000 999.500000 366.350000 ;
      RECT 907.500000 365.650000 949.500000 366.350000 ;
      RECT 857.500000 365.650000 899.500000 366.350000 ;
      RECT 807.500000 365.650000 849.500000 366.350000 ;
      RECT 757.500000 365.650000 799.500000 366.350000 ;
      RECT 707.500000 365.650000 749.500000 366.350000 ;
      RECT 657.500000 365.650000 699.500000 366.350000 ;
      RECT 607.500000 365.650000 649.500000 366.350000 ;
      RECT 557.500000 365.650000 599.500000 366.350000 ;
      RECT 507.500000 365.650000 549.500000 366.350000 ;
      RECT 407.500000 365.650000 449.500000 366.350000 ;
      RECT 357.500000 365.650000 399.500000 366.350000 ;
      RECT 307.500000 365.650000 349.500000 366.350000 ;
      RECT 257.500000 365.650000 299.500000 366.350000 ;
      RECT 207.500000 365.650000 249.500000 366.350000 ;
      RECT 157.500000 365.650000 199.500000 366.350000 ;
      RECT 107.500000 365.650000 149.500000 366.350000 ;
      RECT 57.500000 365.650000 99.500000 366.350000 ;
      RECT 15.500000 365.650000 49.500000 366.350000 ;
      RECT 457.500000 364.605000 499.500000 367.650000 ;
      RECT 416.500000 364.605000 449.500000 365.650000 ;
      RECT 1183.500000 364.350000 1186.000000 367.650000 ;
      RECT 1169.500000 364.350000 1170.500000 365.650000 ;
      RECT 1116.500000 364.350000 1149.500000 365.650000 ;
      RECT 1107.500000 364.350000 1108.500000 365.650000 ;
      RECT 1066.500000 364.350000 1099.500000 365.650000 ;
      RECT 1057.500000 364.350000 1058.500000 365.650000 ;
      RECT 1016.500000 364.350000 1049.500000 365.650000 ;
      RECT 1007.500000 364.350000 1008.500000 365.650000 ;
      RECT 966.500000 364.350000 999.500000 365.650000 ;
      RECT 957.500000 364.350000 958.500000 365.650000 ;
      RECT 916.500000 364.350000 949.500000 365.650000 ;
      RECT 907.500000 364.350000 908.500000 365.650000 ;
      RECT 866.500000 364.350000 899.500000 365.650000 ;
      RECT 857.500000 364.350000 858.500000 365.650000 ;
      RECT 816.500000 364.350000 849.500000 365.650000 ;
      RECT 807.500000 364.350000 808.500000 365.650000 ;
      RECT 766.500000 364.350000 799.500000 365.650000 ;
      RECT 757.500000 364.350000 758.500000 365.650000 ;
      RECT 716.500000 364.350000 749.500000 365.650000 ;
      RECT 707.500000 364.350000 708.500000 365.650000 ;
      RECT 666.500000 364.350000 699.500000 365.650000 ;
      RECT 657.500000 364.350000 658.500000 365.650000 ;
      RECT 616.500000 364.350000 649.500000 365.650000 ;
      RECT 607.500000 364.350000 608.500000 365.650000 ;
      RECT 566.500000 364.350000 599.500000 365.650000 ;
      RECT 557.500000 364.350000 558.500000 365.650000 ;
      RECT 516.500000 364.350000 549.500000 365.650000 ;
      RECT 507.500000 364.350000 508.500000 365.650000 ;
      RECT 416.500000 364.350000 499.500000 364.605000 ;
      RECT 407.500000 364.350000 408.500000 365.650000 ;
      RECT 366.500000 364.350000 399.500000 365.650000 ;
      RECT 357.500000 364.350000 358.500000 365.650000 ;
      RECT 316.500000 364.350000 349.500000 365.650000 ;
      RECT 307.500000 364.350000 308.500000 365.650000 ;
      RECT 266.500000 364.350000 299.500000 365.650000 ;
      RECT 257.500000 364.350000 258.500000 365.650000 ;
      RECT 216.500000 364.350000 249.500000 365.650000 ;
      RECT 207.500000 364.350000 208.500000 365.650000 ;
      RECT 166.500000 364.350000 199.500000 365.650000 ;
      RECT 157.500000 364.350000 158.500000 365.650000 ;
      RECT 116.500000 364.350000 149.500000 365.650000 ;
      RECT 107.500000 364.350000 108.500000 365.650000 ;
      RECT 66.500000 364.350000 99.500000 365.650000 ;
      RECT 57.500000 364.350000 58.500000 365.650000 ;
      RECT 29.500000 364.350000 49.500000 365.650000 ;
      RECT 15.500000 364.350000 16.500000 365.650000 ;
      RECT 0.000000 364.350000 2.500000 367.650000 ;
      RECT 1169.500000 363.650000 1186.000000 364.350000 ;
      RECT 1116.500000 363.650000 1156.500000 364.350000 ;
      RECT 1066.500000 363.650000 1108.500000 364.350000 ;
      RECT 1016.500000 363.650000 1058.500000 364.350000 ;
      RECT 966.500000 363.650000 1008.500000 364.350000 ;
      RECT 916.500000 363.650000 958.500000 364.350000 ;
      RECT 866.500000 363.650000 908.500000 364.350000 ;
      RECT 816.500000 363.650000 858.500000 364.350000 ;
      RECT 766.500000 363.650000 808.500000 364.350000 ;
      RECT 716.500000 363.650000 758.500000 364.350000 ;
      RECT 666.500000 363.650000 708.500000 364.350000 ;
      RECT 616.500000 363.650000 658.500000 364.350000 ;
      RECT 566.500000 363.650000 608.500000 364.350000 ;
      RECT 516.500000 363.650000 558.500000 364.350000 ;
      RECT 416.500000 363.650000 508.500000 364.350000 ;
      RECT 366.500000 363.650000 408.500000 364.350000 ;
      RECT 316.500000 363.650000 358.500000 364.350000 ;
      RECT 266.500000 363.650000 308.500000 364.350000 ;
      RECT 216.500000 363.650000 258.500000 364.350000 ;
      RECT 166.500000 363.650000 208.500000 364.350000 ;
      RECT 116.500000 363.650000 158.500000 364.350000 ;
      RECT 66.500000 363.650000 108.500000 364.350000 ;
      RECT 29.500000 363.650000 58.500000 364.350000 ;
      RECT 0.000000 363.650000 16.500000 364.350000 ;
      RECT 1169.500000 362.350000 1170.500000 363.650000 ;
      RECT 1116.500000 362.350000 1149.500000 363.650000 ;
      RECT 1107.500000 362.350000 1108.500000 363.650000 ;
      RECT 1066.500000 362.350000 1099.500000 363.650000 ;
      RECT 1057.500000 362.350000 1058.500000 363.650000 ;
      RECT 1016.500000 362.350000 1049.500000 363.650000 ;
      RECT 1007.500000 362.350000 1008.500000 363.650000 ;
      RECT 966.500000 362.350000 999.500000 363.650000 ;
      RECT 957.500000 362.350000 958.500000 363.650000 ;
      RECT 916.500000 362.350000 949.500000 363.650000 ;
      RECT 907.500000 362.350000 908.500000 363.650000 ;
      RECT 866.500000 362.350000 899.500000 363.650000 ;
      RECT 857.500000 362.350000 858.500000 363.650000 ;
      RECT 816.500000 362.350000 849.500000 363.650000 ;
      RECT 807.500000 362.350000 808.500000 363.650000 ;
      RECT 766.500000 362.350000 799.500000 363.650000 ;
      RECT 757.500000 362.350000 758.500000 363.650000 ;
      RECT 716.500000 362.350000 749.500000 363.650000 ;
      RECT 707.500000 362.350000 708.500000 363.650000 ;
      RECT 666.500000 362.350000 699.500000 363.650000 ;
      RECT 657.500000 362.350000 658.500000 363.650000 ;
      RECT 616.500000 362.350000 649.500000 363.650000 ;
      RECT 607.500000 362.350000 608.500000 363.650000 ;
      RECT 566.500000 362.350000 599.500000 363.650000 ;
      RECT 557.500000 362.350000 558.500000 363.650000 ;
      RECT 516.500000 362.350000 549.500000 363.650000 ;
      RECT 507.500000 362.350000 508.500000 363.650000 ;
      RECT 416.500000 362.350000 499.500000 363.650000 ;
      RECT 407.500000 362.350000 408.500000 363.650000 ;
      RECT 366.500000 362.350000 399.500000 363.650000 ;
      RECT 357.500000 362.350000 358.500000 363.650000 ;
      RECT 316.500000 362.350000 349.500000 363.650000 ;
      RECT 307.500000 362.350000 308.500000 363.650000 ;
      RECT 266.500000 362.350000 299.500000 363.650000 ;
      RECT 257.500000 362.350000 258.500000 363.650000 ;
      RECT 216.500000 362.350000 249.500000 363.650000 ;
      RECT 207.500000 362.350000 208.500000 363.650000 ;
      RECT 166.500000 362.350000 199.500000 363.650000 ;
      RECT 157.500000 362.350000 158.500000 363.650000 ;
      RECT 116.500000 362.350000 149.500000 363.650000 ;
      RECT 107.500000 362.350000 108.500000 363.650000 ;
      RECT 66.500000 362.350000 99.500000 363.650000 ;
      RECT 57.500000 362.350000 58.500000 363.650000 ;
      RECT 29.500000 362.350000 49.500000 363.650000 ;
      RECT 15.500000 362.350000 16.500000 363.650000 ;
      RECT 1157.500000 361.650000 1170.500000 362.350000 ;
      RECT 1107.500000 361.650000 1149.500000 362.350000 ;
      RECT 1057.500000 361.650000 1099.500000 362.350000 ;
      RECT 1007.500000 361.650000 1049.500000 362.350000 ;
      RECT 957.500000 361.650000 999.500000 362.350000 ;
      RECT 907.500000 361.650000 949.500000 362.350000 ;
      RECT 857.500000 361.650000 899.500000 362.350000 ;
      RECT 807.500000 361.650000 849.500000 362.350000 ;
      RECT 757.500000 361.650000 799.500000 362.350000 ;
      RECT 707.500000 361.650000 749.500000 362.350000 ;
      RECT 657.500000 361.650000 699.500000 362.350000 ;
      RECT 607.500000 361.650000 649.500000 362.350000 ;
      RECT 557.500000 361.650000 599.500000 362.350000 ;
      RECT 507.500000 361.650000 549.500000 362.350000 ;
      RECT 407.500000 361.650000 499.500000 362.350000 ;
      RECT 357.500000 361.650000 399.500000 362.350000 ;
      RECT 307.500000 361.650000 349.500000 362.350000 ;
      RECT 257.500000 361.650000 299.500000 362.350000 ;
      RECT 207.500000 361.650000 249.500000 362.350000 ;
      RECT 157.500000 361.650000 199.500000 362.350000 ;
      RECT 107.500000 361.650000 149.500000 362.350000 ;
      RECT 15.500000 361.650000 49.500000 362.350000 ;
      RECT 1183.500000 360.350000 1186.000000 363.650000 ;
      RECT 1169.500000 360.350000 1170.500000 361.650000 ;
      RECT 1116.500000 360.350000 1149.500000 361.650000 ;
      RECT 1107.500000 360.350000 1108.500000 361.650000 ;
      RECT 1066.500000 360.350000 1099.500000 361.650000 ;
      RECT 1057.500000 360.350000 1058.500000 361.650000 ;
      RECT 1016.500000 360.350000 1049.500000 361.650000 ;
      RECT 1007.500000 360.350000 1008.500000 361.650000 ;
      RECT 966.500000 360.350000 999.500000 361.650000 ;
      RECT 957.500000 360.350000 958.500000 361.650000 ;
      RECT 916.500000 360.350000 949.500000 361.650000 ;
      RECT 907.500000 360.350000 908.500000 361.650000 ;
      RECT 866.500000 360.350000 899.500000 361.650000 ;
      RECT 857.500000 360.350000 858.500000 361.650000 ;
      RECT 816.500000 360.350000 849.500000 361.650000 ;
      RECT 807.500000 360.350000 808.500000 361.650000 ;
      RECT 766.500000 360.350000 799.500000 361.650000 ;
      RECT 757.500000 360.350000 758.500000 361.650000 ;
      RECT 716.500000 360.350000 749.500000 361.650000 ;
      RECT 707.500000 360.350000 708.500000 361.650000 ;
      RECT 666.500000 360.350000 699.500000 361.650000 ;
      RECT 657.500000 360.350000 658.500000 361.650000 ;
      RECT 616.500000 360.350000 649.500000 361.650000 ;
      RECT 607.500000 360.350000 608.500000 361.650000 ;
      RECT 566.500000 360.350000 599.500000 361.650000 ;
      RECT 557.500000 360.350000 558.500000 361.650000 ;
      RECT 516.500000 360.350000 549.500000 361.650000 ;
      RECT 507.500000 360.350000 508.500000 361.650000 ;
      RECT 416.500000 360.350000 499.500000 361.650000 ;
      RECT 407.500000 360.350000 408.500000 361.650000 ;
      RECT 366.500000 360.350000 399.500000 361.650000 ;
      RECT 357.500000 360.350000 358.500000 361.650000 ;
      RECT 316.500000 360.350000 349.500000 361.650000 ;
      RECT 307.500000 360.350000 308.500000 361.650000 ;
      RECT 266.500000 360.350000 299.500000 361.650000 ;
      RECT 257.500000 360.350000 258.500000 361.650000 ;
      RECT 216.500000 360.350000 249.500000 361.650000 ;
      RECT 207.500000 360.350000 208.500000 361.650000 ;
      RECT 166.500000 360.350000 199.500000 361.650000 ;
      RECT 157.500000 360.350000 158.500000 361.650000 ;
      RECT 116.500000 360.350000 149.500000 361.650000 ;
      RECT 107.500000 360.350000 108.500000 361.650000 ;
      RECT 57.500000 360.350000 99.500000 362.350000 ;
      RECT 29.500000 360.350000 49.500000 361.650000 ;
      RECT 15.500000 360.350000 16.500000 361.650000 ;
      RECT 0.000000 360.350000 2.500000 363.650000 ;
      RECT 1169.500000 359.650000 1186.000000 360.350000 ;
      RECT 1116.500000 359.650000 1156.500000 360.350000 ;
      RECT 1066.500000 359.650000 1108.500000 360.350000 ;
      RECT 1016.500000 359.650000 1058.500000 360.350000 ;
      RECT 966.500000 359.650000 1008.500000 360.350000 ;
      RECT 916.500000 359.650000 958.500000 360.350000 ;
      RECT 866.500000 359.650000 908.500000 360.350000 ;
      RECT 816.500000 359.650000 858.500000 360.350000 ;
      RECT 766.500000 359.650000 808.500000 360.350000 ;
      RECT 716.500000 359.650000 758.500000 360.350000 ;
      RECT 666.500000 359.650000 708.500000 360.350000 ;
      RECT 616.500000 359.650000 658.500000 360.350000 ;
      RECT 566.500000 359.650000 608.500000 360.350000 ;
      RECT 516.500000 359.650000 558.500000 360.350000 ;
      RECT 416.500000 359.650000 508.500000 360.350000 ;
      RECT 366.500000 359.650000 408.500000 360.350000 ;
      RECT 316.500000 359.650000 358.500000 360.350000 ;
      RECT 266.500000 359.650000 308.500000 360.350000 ;
      RECT 216.500000 359.650000 258.500000 360.350000 ;
      RECT 166.500000 359.650000 208.500000 360.350000 ;
      RECT 116.500000 359.650000 158.500000 360.350000 ;
      RECT 29.500000 359.650000 108.500000 360.350000 ;
      RECT 0.000000 359.650000 16.500000 360.350000 ;
      RECT 1169.500000 358.350000 1170.500000 359.650000 ;
      RECT 1116.500000 358.350000 1149.500000 359.650000 ;
      RECT 1107.500000 358.350000 1108.500000 359.650000 ;
      RECT 1066.500000 358.350000 1099.500000 359.650000 ;
      RECT 1057.500000 358.350000 1058.500000 359.650000 ;
      RECT 1016.500000 358.350000 1049.500000 359.650000 ;
      RECT 1007.500000 358.350000 1008.500000 359.650000 ;
      RECT 966.500000 358.350000 999.500000 359.650000 ;
      RECT 957.500000 358.350000 958.500000 359.650000 ;
      RECT 916.500000 358.350000 949.500000 359.650000 ;
      RECT 907.500000 358.350000 908.500000 359.650000 ;
      RECT 866.500000 358.350000 899.500000 359.650000 ;
      RECT 857.500000 358.350000 858.500000 359.650000 ;
      RECT 816.500000 358.350000 849.500000 359.650000 ;
      RECT 807.500000 358.350000 808.500000 359.650000 ;
      RECT 766.500000 358.350000 799.500000 359.650000 ;
      RECT 757.500000 358.350000 758.500000 359.650000 ;
      RECT 716.500000 358.350000 749.500000 359.650000 ;
      RECT 707.500000 358.350000 708.500000 359.650000 ;
      RECT 666.500000 358.350000 699.500000 359.650000 ;
      RECT 657.500000 358.350000 658.500000 359.650000 ;
      RECT 616.500000 358.350000 649.500000 359.650000 ;
      RECT 607.500000 358.350000 608.500000 359.650000 ;
      RECT 566.500000 358.350000 599.500000 359.650000 ;
      RECT 557.500000 358.350000 558.500000 359.650000 ;
      RECT 516.500000 358.350000 549.500000 359.650000 ;
      RECT 507.500000 358.350000 508.500000 359.650000 ;
      RECT 416.500000 358.350000 499.500000 359.650000 ;
      RECT 407.500000 358.350000 408.500000 359.650000 ;
      RECT 366.500000 358.350000 399.500000 359.650000 ;
      RECT 357.500000 358.350000 358.500000 359.650000 ;
      RECT 316.500000 358.350000 349.500000 359.650000 ;
      RECT 307.500000 358.350000 308.500000 359.650000 ;
      RECT 266.500000 358.350000 299.500000 359.650000 ;
      RECT 257.500000 358.350000 258.500000 359.650000 ;
      RECT 216.500000 358.350000 249.500000 359.650000 ;
      RECT 207.500000 358.350000 208.500000 359.650000 ;
      RECT 166.500000 358.350000 199.500000 359.650000 ;
      RECT 157.500000 358.350000 158.500000 359.650000 ;
      RECT 116.500000 358.350000 149.500000 359.650000 ;
      RECT 107.500000 358.350000 108.500000 359.650000 ;
      RECT 29.500000 358.350000 99.500000 359.650000 ;
      RECT 15.500000 358.350000 16.500000 359.650000 ;
      RECT 1157.500000 357.650000 1170.500000 358.350000 ;
      RECT 1107.500000 357.650000 1149.500000 358.350000 ;
      RECT 1057.500000 357.650000 1099.500000 358.350000 ;
      RECT 1007.500000 357.650000 1049.500000 358.350000 ;
      RECT 957.500000 357.650000 999.500000 358.350000 ;
      RECT 907.500000 357.650000 949.500000 358.350000 ;
      RECT 857.500000 357.650000 899.500000 358.350000 ;
      RECT 807.500000 357.650000 849.500000 358.350000 ;
      RECT 757.500000 357.650000 799.500000 358.350000 ;
      RECT 707.500000 357.650000 749.500000 358.350000 ;
      RECT 657.500000 357.650000 699.500000 358.350000 ;
      RECT 607.500000 357.650000 649.500000 358.350000 ;
      RECT 557.500000 357.650000 599.500000 358.350000 ;
      RECT 507.500000 357.650000 549.500000 358.350000 ;
      RECT 407.500000 357.650000 499.500000 358.350000 ;
      RECT 357.500000 357.650000 399.500000 358.350000 ;
      RECT 307.500000 357.650000 349.500000 358.350000 ;
      RECT 257.500000 357.650000 299.500000 358.350000 ;
      RECT 207.500000 357.650000 249.500000 358.350000 ;
      RECT 157.500000 357.650000 199.500000 358.350000 ;
      RECT 107.500000 357.650000 149.500000 358.350000 ;
      RECT 15.500000 357.650000 99.500000 358.350000 ;
      RECT 1183.500000 356.350000 1186.000000 359.650000 ;
      RECT 1169.500000 356.350000 1170.500000 357.650000 ;
      RECT 1116.500000 356.350000 1149.500000 357.650000 ;
      RECT 1107.500000 356.350000 1108.500000 357.650000 ;
      RECT 1066.500000 356.350000 1099.500000 357.650000 ;
      RECT 1057.500000 356.350000 1058.500000 357.650000 ;
      RECT 1016.500000 356.350000 1049.500000 357.650000 ;
      RECT 1007.500000 356.350000 1008.500000 357.650000 ;
      RECT 966.500000 356.350000 999.500000 357.650000 ;
      RECT 957.500000 356.350000 958.500000 357.650000 ;
      RECT 916.500000 356.350000 949.500000 357.650000 ;
      RECT 907.500000 356.350000 908.500000 357.650000 ;
      RECT 866.500000 356.350000 899.500000 357.650000 ;
      RECT 857.500000 356.350000 858.500000 357.650000 ;
      RECT 816.500000 356.350000 849.500000 357.650000 ;
      RECT 807.500000 356.350000 808.500000 357.650000 ;
      RECT 766.500000 356.350000 799.500000 357.650000 ;
      RECT 757.500000 356.350000 758.500000 357.650000 ;
      RECT 716.500000 356.350000 749.500000 357.650000 ;
      RECT 707.500000 356.350000 708.500000 357.650000 ;
      RECT 666.500000 356.350000 699.500000 357.650000 ;
      RECT 657.500000 356.350000 658.500000 357.650000 ;
      RECT 616.500000 356.350000 649.500000 357.650000 ;
      RECT 607.500000 356.350000 608.500000 357.650000 ;
      RECT 566.500000 356.350000 599.500000 357.650000 ;
      RECT 557.500000 356.350000 558.500000 357.650000 ;
      RECT 516.500000 356.350000 549.500000 357.650000 ;
      RECT 507.500000 356.350000 508.500000 357.650000 ;
      RECT 416.500000 356.350000 499.500000 357.650000 ;
      RECT 407.500000 356.350000 408.500000 357.650000 ;
      RECT 366.500000 356.350000 399.500000 357.650000 ;
      RECT 357.500000 356.350000 358.500000 357.650000 ;
      RECT 316.500000 356.350000 349.500000 357.650000 ;
      RECT 307.500000 356.350000 308.500000 357.650000 ;
      RECT 266.500000 356.350000 299.500000 357.650000 ;
      RECT 257.500000 356.350000 258.500000 357.650000 ;
      RECT 216.500000 356.350000 249.500000 357.650000 ;
      RECT 207.500000 356.350000 208.500000 357.650000 ;
      RECT 166.500000 356.350000 199.500000 357.650000 ;
      RECT 157.500000 356.350000 158.500000 357.650000 ;
      RECT 116.500000 356.350000 149.500000 357.650000 ;
      RECT 107.500000 356.350000 108.500000 357.650000 ;
      RECT 29.500000 356.350000 99.500000 357.650000 ;
      RECT 15.500000 356.350000 16.500000 357.650000 ;
      RECT 0.000000 356.350000 2.500000 359.650000 ;
      RECT 29.500000 356.245000 108.500000 356.350000 ;
      RECT 1169.500000 355.650000 1186.000000 356.350000 ;
      RECT 1116.500000 355.650000 1156.500000 356.350000 ;
      RECT 1066.500000 355.650000 1108.500000 356.350000 ;
      RECT 1016.500000 355.650000 1058.500000 356.350000 ;
      RECT 966.500000 355.650000 1008.500000 356.350000 ;
      RECT 916.500000 355.650000 958.500000 356.350000 ;
      RECT 866.500000 355.650000 908.500000 356.350000 ;
      RECT 816.500000 355.650000 858.500000 356.350000 ;
      RECT 766.500000 355.650000 808.500000 356.350000 ;
      RECT 716.500000 355.650000 758.500000 356.350000 ;
      RECT 666.500000 355.650000 708.500000 356.350000 ;
      RECT 616.500000 355.650000 658.500000 356.350000 ;
      RECT 566.500000 355.650000 608.500000 356.350000 ;
      RECT 516.500000 355.650000 558.500000 356.350000 ;
      RECT 416.500000 355.650000 508.500000 356.350000 ;
      RECT 366.500000 355.650000 408.500000 356.350000 ;
      RECT 316.500000 355.650000 358.500000 356.350000 ;
      RECT 266.500000 355.650000 308.500000 356.350000 ;
      RECT 216.500000 355.650000 258.500000 356.350000 ;
      RECT 166.500000 355.650000 208.500000 356.350000 ;
      RECT 116.500000 355.650000 158.500000 356.350000 ;
      RECT 57.500000 355.650000 108.500000 356.245000 ;
      RECT 0.000000 355.650000 16.500000 356.350000 ;
      RECT 1169.500000 354.350000 1170.500000 355.650000 ;
      RECT 1116.500000 354.350000 1149.500000 355.650000 ;
      RECT 1107.500000 354.350000 1108.500000 355.650000 ;
      RECT 1066.500000 354.350000 1099.500000 355.650000 ;
      RECT 1057.500000 354.350000 1058.500000 355.650000 ;
      RECT 1016.500000 354.350000 1049.500000 355.650000 ;
      RECT 1007.500000 354.350000 1008.500000 355.650000 ;
      RECT 966.500000 354.350000 999.500000 355.650000 ;
      RECT 957.500000 354.350000 958.500000 355.650000 ;
      RECT 916.500000 354.350000 949.500000 355.650000 ;
      RECT 907.500000 354.350000 908.500000 355.650000 ;
      RECT 866.500000 354.350000 899.500000 355.650000 ;
      RECT 857.500000 354.350000 858.500000 355.650000 ;
      RECT 816.500000 354.350000 849.500000 355.650000 ;
      RECT 807.500000 354.350000 808.500000 355.650000 ;
      RECT 766.500000 354.350000 799.500000 355.650000 ;
      RECT 757.500000 354.350000 758.500000 355.650000 ;
      RECT 716.500000 354.350000 749.500000 355.650000 ;
      RECT 707.500000 354.350000 708.500000 355.650000 ;
      RECT 666.500000 354.350000 699.500000 355.650000 ;
      RECT 657.500000 354.350000 658.500000 355.650000 ;
      RECT 616.500000 354.350000 649.500000 355.650000 ;
      RECT 607.500000 354.350000 608.500000 355.650000 ;
      RECT 566.500000 354.350000 599.500000 355.650000 ;
      RECT 557.500000 354.350000 558.500000 355.650000 ;
      RECT 516.500000 354.350000 549.500000 355.650000 ;
      RECT 507.500000 354.350000 508.500000 355.650000 ;
      RECT 416.500000 354.350000 499.500000 355.650000 ;
      RECT 407.500000 354.350000 408.500000 355.650000 ;
      RECT 366.500000 354.350000 399.500000 355.650000 ;
      RECT 357.500000 354.350000 358.500000 355.650000 ;
      RECT 316.500000 354.350000 349.500000 355.650000 ;
      RECT 307.500000 354.350000 308.500000 355.650000 ;
      RECT 266.500000 354.350000 299.500000 355.650000 ;
      RECT 257.500000 354.350000 258.500000 355.650000 ;
      RECT 216.500000 354.350000 249.500000 355.650000 ;
      RECT 207.500000 354.350000 208.500000 355.650000 ;
      RECT 166.500000 354.350000 199.500000 355.650000 ;
      RECT 157.500000 354.350000 158.500000 355.650000 ;
      RECT 116.500000 354.350000 149.500000 355.650000 ;
      RECT 107.500000 354.350000 108.500000 355.650000 ;
      RECT 29.500000 354.350000 49.500000 356.245000 ;
      RECT 15.500000 354.350000 16.500000 355.650000 ;
      RECT 57.500000 354.245000 99.500000 355.650000 ;
      RECT 407.500000 353.730000 499.500000 354.350000 ;
      RECT 1157.500000 353.650000 1170.500000 354.350000 ;
      RECT 1107.500000 353.650000 1149.500000 354.350000 ;
      RECT 1057.500000 353.650000 1099.500000 354.350000 ;
      RECT 1007.500000 353.650000 1049.500000 354.350000 ;
      RECT 957.500000 353.650000 999.500000 354.350000 ;
      RECT 907.500000 353.650000 949.500000 354.350000 ;
      RECT 857.500000 353.650000 899.500000 354.350000 ;
      RECT 807.500000 353.650000 849.500000 354.350000 ;
      RECT 757.500000 353.650000 799.500000 354.350000 ;
      RECT 707.500000 353.650000 749.500000 354.350000 ;
      RECT 657.500000 353.650000 699.500000 354.350000 ;
      RECT 607.500000 353.650000 649.500000 354.350000 ;
      RECT 557.500000 353.650000 599.500000 354.350000 ;
      RECT 507.500000 353.650000 549.500000 354.350000 ;
      RECT 407.500000 353.650000 458.500000 353.730000 ;
      RECT 357.500000 353.650000 399.500000 354.350000 ;
      RECT 307.500000 353.650000 349.500000 354.350000 ;
      RECT 257.500000 353.650000 299.500000 354.350000 ;
      RECT 207.500000 353.650000 249.500000 354.350000 ;
      RECT 157.500000 353.650000 199.500000 354.350000 ;
      RECT 107.500000 353.650000 149.500000 354.350000 ;
      RECT 15.500000 353.650000 49.500000 354.350000 ;
      RECT 57.500000 352.945000 58.500000 354.245000 ;
      RECT 29.500000 352.945000 49.500000 353.650000 ;
      RECT 1183.500000 352.350000 1186.000000 355.650000 ;
      RECT 1169.500000 352.350000 1170.500000 353.650000 ;
      RECT 1116.500000 352.350000 1149.500000 353.650000 ;
      RECT 1107.500000 352.350000 1108.500000 353.650000 ;
      RECT 1066.500000 352.350000 1099.500000 353.650000 ;
      RECT 1057.500000 352.350000 1058.500000 353.650000 ;
      RECT 1016.500000 352.350000 1049.500000 353.650000 ;
      RECT 1007.500000 352.350000 1008.500000 353.650000 ;
      RECT 966.500000 352.350000 999.500000 353.650000 ;
      RECT 957.500000 352.350000 958.500000 353.650000 ;
      RECT 916.500000 352.350000 949.500000 353.650000 ;
      RECT 907.500000 352.350000 908.500000 353.650000 ;
      RECT 866.500000 352.350000 899.500000 353.650000 ;
      RECT 857.500000 352.350000 858.500000 353.650000 ;
      RECT 816.500000 352.350000 849.500000 353.650000 ;
      RECT 807.500000 352.350000 808.500000 353.650000 ;
      RECT 766.500000 352.350000 799.500000 353.650000 ;
      RECT 757.500000 352.350000 758.500000 353.650000 ;
      RECT 716.500000 352.350000 749.500000 353.650000 ;
      RECT 707.500000 352.350000 708.500000 353.650000 ;
      RECT 666.500000 352.350000 699.500000 353.650000 ;
      RECT 657.500000 352.350000 658.500000 353.650000 ;
      RECT 616.500000 352.350000 649.500000 353.650000 ;
      RECT 607.500000 352.350000 608.500000 353.650000 ;
      RECT 566.500000 352.350000 599.500000 353.650000 ;
      RECT 557.500000 352.350000 558.500000 353.650000 ;
      RECT 516.500000 352.350000 549.500000 353.650000 ;
      RECT 507.500000 352.350000 508.500000 353.650000 ;
      RECT 466.500000 352.350000 499.500000 353.730000 ;
      RECT 407.500000 352.350000 408.500000 353.650000 ;
      RECT 366.500000 352.350000 399.500000 353.650000 ;
      RECT 357.500000 352.350000 358.500000 353.650000 ;
      RECT 316.500000 352.350000 349.500000 353.650000 ;
      RECT 307.500000 352.350000 308.500000 353.650000 ;
      RECT 266.500000 352.350000 299.500000 353.650000 ;
      RECT 257.500000 352.350000 258.500000 353.650000 ;
      RECT 216.500000 352.350000 249.500000 353.650000 ;
      RECT 207.500000 352.350000 208.500000 353.650000 ;
      RECT 166.500000 352.350000 199.500000 353.650000 ;
      RECT 157.500000 352.350000 158.500000 353.650000 ;
      RECT 116.500000 352.350000 149.500000 353.650000 ;
      RECT 107.500000 352.350000 108.500000 353.650000 ;
      RECT 65.580000 352.350000 99.500000 354.245000 ;
      RECT 15.500000 352.350000 16.500000 353.650000 ;
      RECT 0.000000 352.350000 2.500000 355.650000 ;
      RECT 1169.500000 351.650000 1186.000000 352.350000 ;
      RECT 1116.500000 351.650000 1156.500000 352.350000 ;
      RECT 1066.500000 351.650000 1108.500000 352.350000 ;
      RECT 1016.500000 351.650000 1058.500000 352.350000 ;
      RECT 966.500000 351.650000 1008.500000 352.350000 ;
      RECT 916.500000 351.650000 958.500000 352.350000 ;
      RECT 866.500000 351.650000 908.500000 352.350000 ;
      RECT 816.500000 351.650000 858.500000 352.350000 ;
      RECT 766.500000 351.650000 808.500000 352.350000 ;
      RECT 716.500000 351.650000 758.500000 352.350000 ;
      RECT 666.500000 351.650000 708.500000 352.350000 ;
      RECT 616.500000 351.650000 658.500000 352.350000 ;
      RECT 566.500000 351.650000 608.500000 352.350000 ;
      RECT 516.500000 351.650000 558.500000 352.350000 ;
      RECT 466.500000 351.650000 508.500000 352.350000 ;
      RECT 366.500000 351.650000 408.500000 352.350000 ;
      RECT 316.500000 351.650000 358.500000 352.350000 ;
      RECT 266.500000 351.650000 308.500000 352.350000 ;
      RECT 216.500000 351.650000 258.500000 352.350000 ;
      RECT 166.500000 351.650000 208.500000 352.350000 ;
      RECT 116.500000 351.650000 158.500000 352.350000 ;
      RECT 65.580000 351.650000 108.500000 352.350000 ;
      RECT 0.000000 351.650000 16.500000 352.350000 ;
      RECT 65.580000 350.945000 99.500000 351.650000 ;
      RECT 29.500000 350.945000 58.500000 352.945000 ;
      RECT 1169.500000 350.350000 1170.500000 351.650000 ;
      RECT 1116.500000 350.350000 1149.500000 351.650000 ;
      RECT 1107.500000 350.350000 1108.500000 351.650000 ;
      RECT 1066.500000 350.350000 1099.500000 351.650000 ;
      RECT 1057.500000 350.350000 1058.500000 351.650000 ;
      RECT 1016.500000 350.350000 1049.500000 351.650000 ;
      RECT 1007.500000 350.350000 1008.500000 351.650000 ;
      RECT 966.500000 350.350000 999.500000 351.650000 ;
      RECT 957.500000 350.350000 958.500000 351.650000 ;
      RECT 916.500000 350.350000 949.500000 351.650000 ;
      RECT 907.500000 350.350000 908.500000 351.650000 ;
      RECT 866.500000 350.350000 899.500000 351.650000 ;
      RECT 857.500000 350.350000 858.500000 351.650000 ;
      RECT 816.500000 350.350000 849.500000 351.650000 ;
      RECT 807.500000 350.350000 808.500000 351.650000 ;
      RECT 766.500000 350.350000 799.500000 351.650000 ;
      RECT 757.500000 350.350000 758.500000 351.650000 ;
      RECT 716.500000 350.350000 749.500000 351.650000 ;
      RECT 707.500000 350.350000 708.500000 351.650000 ;
      RECT 666.500000 350.350000 699.500000 351.650000 ;
      RECT 657.500000 350.350000 658.500000 351.650000 ;
      RECT 616.500000 350.350000 649.500000 351.650000 ;
      RECT 607.500000 350.350000 608.500000 351.650000 ;
      RECT 566.500000 350.350000 599.500000 351.650000 ;
      RECT 557.500000 350.350000 558.500000 351.650000 ;
      RECT 516.500000 350.350000 549.500000 351.650000 ;
      RECT 507.500000 350.350000 508.500000 351.650000 ;
      RECT 416.500000 350.350000 458.500000 353.650000 ;
      RECT 407.500000 350.350000 408.500000 351.650000 ;
      RECT 366.500000 350.350000 399.500000 351.650000 ;
      RECT 357.500000 350.350000 358.500000 351.650000 ;
      RECT 316.500000 350.350000 349.500000 351.650000 ;
      RECT 307.500000 350.350000 308.500000 351.650000 ;
      RECT 266.500000 350.350000 299.500000 351.650000 ;
      RECT 257.500000 350.350000 258.500000 351.650000 ;
      RECT 216.500000 350.350000 249.500000 351.650000 ;
      RECT 207.500000 350.350000 208.500000 351.650000 ;
      RECT 166.500000 350.350000 199.500000 351.650000 ;
      RECT 157.500000 350.350000 158.500000 351.650000 ;
      RECT 116.500000 350.350000 149.500000 351.650000 ;
      RECT 107.500000 350.350000 108.500000 351.650000 ;
      RECT 29.500000 350.350000 99.500000 350.945000 ;
      RECT 15.500000 350.350000 16.500000 351.650000 ;
      RECT 466.500000 349.730000 499.500000 351.650000 ;
      RECT 407.500000 349.730000 458.500000 350.350000 ;
      RECT 1157.500000 349.650000 1170.500000 350.350000 ;
      RECT 1107.500000 349.650000 1149.500000 350.350000 ;
      RECT 1057.500000 349.650000 1099.500000 350.350000 ;
      RECT 1007.500000 349.650000 1049.500000 350.350000 ;
      RECT 957.500000 349.650000 999.500000 350.350000 ;
      RECT 907.500000 349.650000 949.500000 350.350000 ;
      RECT 857.500000 349.650000 899.500000 350.350000 ;
      RECT 807.500000 349.650000 849.500000 350.350000 ;
      RECT 757.500000 349.650000 799.500000 350.350000 ;
      RECT 707.500000 349.650000 749.500000 350.350000 ;
      RECT 657.500000 349.650000 699.500000 350.350000 ;
      RECT 607.500000 349.650000 649.500000 350.350000 ;
      RECT 557.500000 349.650000 599.500000 350.350000 ;
      RECT 507.500000 349.650000 549.500000 350.350000 ;
      RECT 407.500000 349.650000 499.500000 349.730000 ;
      RECT 357.500000 349.650000 399.500000 350.350000 ;
      RECT 307.500000 349.650000 349.500000 350.350000 ;
      RECT 257.500000 349.650000 299.500000 350.350000 ;
      RECT 207.500000 349.650000 249.500000 350.350000 ;
      RECT 157.500000 349.650000 199.500000 350.350000 ;
      RECT 107.500000 349.650000 149.500000 350.350000 ;
      RECT 15.500000 349.650000 99.500000 350.350000 ;
      RECT 1183.500000 348.350000 1186.000000 351.650000 ;
      RECT 1169.500000 348.350000 1170.500000 349.650000 ;
      RECT 1116.500000 348.350000 1149.500000 349.650000 ;
      RECT 1107.500000 348.350000 1108.500000 349.650000 ;
      RECT 1066.500000 348.350000 1099.500000 349.650000 ;
      RECT 1057.500000 348.350000 1058.500000 349.650000 ;
      RECT 1016.500000 348.350000 1049.500000 349.650000 ;
      RECT 1007.500000 348.350000 1008.500000 349.650000 ;
      RECT 966.500000 348.350000 999.500000 349.650000 ;
      RECT 957.500000 348.350000 958.500000 349.650000 ;
      RECT 916.500000 348.350000 949.500000 349.650000 ;
      RECT 907.500000 348.350000 908.500000 349.650000 ;
      RECT 866.500000 348.350000 899.500000 349.650000 ;
      RECT 857.500000 348.350000 858.500000 349.650000 ;
      RECT 816.500000 348.350000 849.500000 349.650000 ;
      RECT 807.500000 348.350000 808.500000 349.650000 ;
      RECT 766.500000 348.350000 799.500000 349.650000 ;
      RECT 757.500000 348.350000 758.500000 349.650000 ;
      RECT 716.500000 348.350000 749.500000 349.650000 ;
      RECT 707.500000 348.350000 708.500000 349.650000 ;
      RECT 666.500000 348.350000 699.500000 349.650000 ;
      RECT 657.500000 348.350000 658.500000 349.650000 ;
      RECT 616.500000 348.350000 649.500000 349.650000 ;
      RECT 607.500000 348.350000 608.500000 349.650000 ;
      RECT 566.500000 348.350000 599.500000 349.650000 ;
      RECT 557.500000 348.350000 558.500000 349.650000 ;
      RECT 516.500000 348.350000 549.500000 349.650000 ;
      RECT 507.500000 348.350000 508.500000 349.650000 ;
      RECT 466.500000 348.350000 499.500000 349.650000 ;
      RECT 407.500000 348.350000 408.500000 349.650000 ;
      RECT 366.500000 348.350000 399.500000 349.650000 ;
      RECT 357.500000 348.350000 358.500000 349.650000 ;
      RECT 316.500000 348.350000 349.500000 349.650000 ;
      RECT 307.500000 348.350000 308.500000 349.650000 ;
      RECT 266.500000 348.350000 299.500000 349.650000 ;
      RECT 257.500000 348.350000 258.500000 349.650000 ;
      RECT 216.500000 348.350000 249.500000 349.650000 ;
      RECT 207.500000 348.350000 208.500000 349.650000 ;
      RECT 166.500000 348.350000 199.500000 349.650000 ;
      RECT 157.500000 348.350000 158.500000 349.650000 ;
      RECT 116.500000 348.350000 149.500000 349.650000 ;
      RECT 107.500000 348.350000 108.500000 349.650000 ;
      RECT 66.500000 348.350000 99.500000 349.650000 ;
      RECT 15.500000 348.350000 16.500000 349.650000 ;
      RECT 0.000000 348.350000 2.500000 351.650000 ;
      RECT 1169.500000 347.650000 1186.000000 348.350000 ;
      RECT 1116.500000 347.650000 1156.500000 348.350000 ;
      RECT 1066.500000 347.650000 1108.500000 348.350000 ;
      RECT 1016.500000 347.650000 1058.500000 348.350000 ;
      RECT 966.500000 347.650000 1008.500000 348.350000 ;
      RECT 916.500000 347.650000 958.500000 348.350000 ;
      RECT 866.500000 347.650000 908.500000 348.350000 ;
      RECT 816.500000 347.650000 858.500000 348.350000 ;
      RECT 766.500000 347.650000 808.500000 348.350000 ;
      RECT 716.500000 347.650000 758.500000 348.350000 ;
      RECT 666.500000 347.650000 708.500000 348.350000 ;
      RECT 616.500000 347.650000 658.500000 348.350000 ;
      RECT 566.500000 347.650000 608.500000 348.350000 ;
      RECT 516.500000 347.650000 558.500000 348.350000 ;
      RECT 466.500000 347.650000 508.500000 348.350000 ;
      RECT 416.500000 347.650000 458.500000 349.650000 ;
      RECT 366.500000 347.650000 408.500000 348.350000 ;
      RECT 316.500000 347.650000 358.500000 348.350000 ;
      RECT 266.500000 347.650000 308.500000 348.350000 ;
      RECT 216.500000 347.650000 258.500000 348.350000 ;
      RECT 166.500000 347.650000 208.500000 348.350000 ;
      RECT 116.500000 347.650000 158.500000 348.350000 ;
      RECT 66.500000 347.650000 108.500000 348.350000 ;
      RECT 29.500000 347.650000 58.500000 349.650000 ;
      RECT 0.000000 347.650000 16.500000 348.350000 ;
      RECT 1169.500000 346.350000 1170.500000 347.650000 ;
      RECT 1116.500000 346.350000 1149.500000 347.650000 ;
      RECT 1107.500000 346.350000 1108.500000 347.650000 ;
      RECT 1066.500000 346.350000 1099.500000 347.650000 ;
      RECT 1057.500000 346.350000 1058.500000 347.650000 ;
      RECT 1016.500000 346.350000 1049.500000 347.650000 ;
      RECT 1007.500000 346.350000 1008.500000 347.650000 ;
      RECT 966.500000 346.350000 999.500000 347.650000 ;
      RECT 957.500000 346.350000 958.500000 347.650000 ;
      RECT 916.500000 346.350000 949.500000 347.650000 ;
      RECT 907.500000 346.350000 908.500000 347.650000 ;
      RECT 866.500000 346.350000 899.500000 347.650000 ;
      RECT 857.500000 346.350000 858.500000 347.650000 ;
      RECT 816.500000 346.350000 849.500000 347.650000 ;
      RECT 807.500000 346.350000 808.500000 347.650000 ;
      RECT 766.500000 346.350000 799.500000 347.650000 ;
      RECT 757.500000 346.350000 758.500000 347.650000 ;
      RECT 716.500000 346.350000 749.500000 347.650000 ;
      RECT 707.500000 346.350000 708.500000 347.650000 ;
      RECT 666.500000 346.350000 699.500000 347.650000 ;
      RECT 657.500000 346.350000 658.500000 347.650000 ;
      RECT 616.500000 346.350000 649.500000 347.650000 ;
      RECT 607.500000 346.350000 608.500000 347.650000 ;
      RECT 566.500000 346.350000 599.500000 347.650000 ;
      RECT 557.500000 346.350000 558.500000 347.650000 ;
      RECT 516.500000 346.350000 549.500000 347.650000 ;
      RECT 507.500000 346.350000 508.500000 347.650000 ;
      RECT 466.500000 346.350000 499.500000 347.650000 ;
      RECT 457.500000 346.350000 458.500000 347.650000 ;
      RECT 416.500000 346.350000 449.500000 347.650000 ;
      RECT 407.500000 346.350000 408.500000 347.650000 ;
      RECT 366.500000 346.350000 399.500000 347.650000 ;
      RECT 357.500000 346.350000 358.500000 347.650000 ;
      RECT 316.500000 346.350000 349.500000 347.650000 ;
      RECT 307.500000 346.350000 308.500000 347.650000 ;
      RECT 266.500000 346.350000 299.500000 347.650000 ;
      RECT 257.500000 346.350000 258.500000 347.650000 ;
      RECT 216.500000 346.350000 249.500000 347.650000 ;
      RECT 207.500000 346.350000 208.500000 347.650000 ;
      RECT 166.500000 346.350000 199.500000 347.650000 ;
      RECT 157.500000 346.350000 158.500000 347.650000 ;
      RECT 116.500000 346.350000 149.500000 347.650000 ;
      RECT 107.500000 346.350000 108.500000 347.650000 ;
      RECT 66.500000 346.350000 99.500000 347.650000 ;
      RECT 57.500000 346.350000 58.500000 347.650000 ;
      RECT 29.500000 346.350000 49.500000 347.650000 ;
      RECT 15.500000 346.350000 16.500000 347.650000 ;
      RECT 1157.500000 345.650000 1170.500000 346.350000 ;
      RECT 1107.500000 345.650000 1149.500000 346.350000 ;
      RECT 1057.500000 345.650000 1099.500000 346.350000 ;
      RECT 1007.500000 345.650000 1049.500000 346.350000 ;
      RECT 957.500000 345.650000 999.500000 346.350000 ;
      RECT 907.500000 345.650000 949.500000 346.350000 ;
      RECT 857.500000 345.650000 899.500000 346.350000 ;
      RECT 807.500000 345.650000 849.500000 346.350000 ;
      RECT 757.500000 345.650000 799.500000 346.350000 ;
      RECT 707.500000 345.650000 749.500000 346.350000 ;
      RECT 657.500000 345.650000 699.500000 346.350000 ;
      RECT 607.500000 345.650000 649.500000 346.350000 ;
      RECT 557.500000 345.650000 599.500000 346.350000 ;
      RECT 507.500000 345.650000 549.500000 346.350000 ;
      RECT 457.500000 345.650000 499.500000 346.350000 ;
      RECT 407.500000 345.650000 449.500000 346.350000 ;
      RECT 357.500000 345.650000 399.500000 346.350000 ;
      RECT 307.500000 345.650000 349.500000 346.350000 ;
      RECT 257.500000 345.650000 299.500000 346.350000 ;
      RECT 207.500000 345.650000 249.500000 346.350000 ;
      RECT 157.500000 345.650000 199.500000 346.350000 ;
      RECT 107.500000 345.650000 149.500000 346.350000 ;
      RECT 57.500000 345.650000 99.500000 346.350000 ;
      RECT 15.500000 345.650000 49.500000 346.350000 ;
      RECT 1183.500000 344.350000 1186.000000 347.650000 ;
      RECT 1169.500000 344.350000 1170.500000 345.650000 ;
      RECT 1116.500000 344.350000 1149.500000 345.650000 ;
      RECT 1107.500000 344.350000 1108.500000 345.650000 ;
      RECT 1066.500000 344.350000 1099.500000 345.650000 ;
      RECT 1057.500000 344.350000 1058.500000 345.650000 ;
      RECT 1016.500000 344.350000 1049.500000 345.650000 ;
      RECT 1007.500000 344.350000 1008.500000 345.650000 ;
      RECT 966.500000 344.350000 999.500000 345.650000 ;
      RECT 957.500000 344.350000 958.500000 345.650000 ;
      RECT 916.500000 344.350000 949.500000 345.650000 ;
      RECT 907.500000 344.350000 908.500000 345.650000 ;
      RECT 866.500000 344.350000 899.500000 345.650000 ;
      RECT 857.500000 344.350000 858.500000 345.650000 ;
      RECT 816.500000 344.350000 849.500000 345.650000 ;
      RECT 807.500000 344.350000 808.500000 345.650000 ;
      RECT 766.500000 344.350000 799.500000 345.650000 ;
      RECT 757.500000 344.350000 758.500000 345.650000 ;
      RECT 716.500000 344.350000 749.500000 345.650000 ;
      RECT 707.500000 344.350000 708.500000 345.650000 ;
      RECT 666.500000 344.350000 699.500000 345.650000 ;
      RECT 657.500000 344.350000 658.500000 345.650000 ;
      RECT 616.500000 344.350000 649.500000 345.650000 ;
      RECT 607.500000 344.350000 608.500000 345.650000 ;
      RECT 566.500000 344.350000 599.500000 345.650000 ;
      RECT 557.500000 344.350000 558.500000 345.650000 ;
      RECT 516.500000 344.350000 549.500000 345.650000 ;
      RECT 507.500000 344.350000 508.500000 345.650000 ;
      RECT 466.500000 344.350000 499.500000 345.650000 ;
      RECT 457.500000 344.350000 458.500000 345.650000 ;
      RECT 416.500000 344.350000 449.500000 345.650000 ;
      RECT 407.500000 344.350000 408.500000 345.650000 ;
      RECT 366.500000 344.350000 399.500000 345.650000 ;
      RECT 357.500000 344.350000 358.500000 345.650000 ;
      RECT 316.500000 344.350000 349.500000 345.650000 ;
      RECT 307.500000 344.350000 308.500000 345.650000 ;
      RECT 266.500000 344.350000 299.500000 345.650000 ;
      RECT 257.500000 344.350000 258.500000 345.650000 ;
      RECT 216.500000 344.350000 249.500000 345.650000 ;
      RECT 207.500000 344.350000 208.500000 345.650000 ;
      RECT 166.500000 344.350000 199.500000 345.650000 ;
      RECT 157.500000 344.350000 158.500000 345.650000 ;
      RECT 116.500000 344.350000 149.500000 345.650000 ;
      RECT 107.500000 344.350000 108.500000 345.650000 ;
      RECT 66.500000 344.350000 99.500000 345.650000 ;
      RECT 57.500000 344.350000 58.500000 345.650000 ;
      RECT 29.500000 344.350000 49.500000 345.650000 ;
      RECT 15.500000 344.350000 16.500000 345.650000 ;
      RECT 0.000000 344.350000 2.500000 347.650000 ;
      RECT 1169.500000 343.650000 1186.000000 344.350000 ;
      RECT 1116.500000 343.650000 1156.500000 344.350000 ;
      RECT 1066.500000 343.650000 1108.500000 344.350000 ;
      RECT 1016.500000 343.650000 1058.500000 344.350000 ;
      RECT 966.500000 343.650000 1008.500000 344.350000 ;
      RECT 916.500000 343.650000 958.500000 344.350000 ;
      RECT 866.500000 343.650000 908.500000 344.350000 ;
      RECT 816.500000 343.650000 858.500000 344.350000 ;
      RECT 766.500000 343.650000 808.500000 344.350000 ;
      RECT 716.500000 343.650000 758.500000 344.350000 ;
      RECT 666.500000 343.650000 708.500000 344.350000 ;
      RECT 616.500000 343.650000 658.500000 344.350000 ;
      RECT 566.500000 343.650000 608.500000 344.350000 ;
      RECT 516.500000 343.650000 558.500000 344.350000 ;
      RECT 466.500000 343.650000 508.500000 344.350000 ;
      RECT 416.500000 343.650000 458.500000 344.350000 ;
      RECT 366.500000 343.650000 408.500000 344.350000 ;
      RECT 316.500000 343.650000 358.500000 344.350000 ;
      RECT 266.500000 343.650000 308.500000 344.350000 ;
      RECT 216.500000 343.650000 258.500000 344.350000 ;
      RECT 166.500000 343.650000 208.500000 344.350000 ;
      RECT 116.500000 343.650000 158.500000 344.350000 ;
      RECT 66.500000 343.650000 108.500000 344.350000 ;
      RECT 29.500000 343.650000 58.500000 344.350000 ;
      RECT 0.000000 343.650000 16.500000 344.350000 ;
      RECT 1169.500000 342.350000 1170.500000 343.650000 ;
      RECT 1116.500000 342.350000 1149.500000 343.650000 ;
      RECT 1107.500000 342.350000 1108.500000 343.650000 ;
      RECT 1066.500000 342.350000 1099.500000 343.650000 ;
      RECT 1057.500000 342.350000 1058.500000 343.650000 ;
      RECT 1016.500000 342.350000 1049.500000 343.650000 ;
      RECT 1007.500000 342.350000 1008.500000 343.650000 ;
      RECT 966.500000 342.350000 999.500000 343.650000 ;
      RECT 957.500000 342.350000 958.500000 343.650000 ;
      RECT 916.500000 342.350000 949.500000 343.650000 ;
      RECT 907.500000 342.350000 908.500000 343.650000 ;
      RECT 866.500000 342.350000 899.500000 343.650000 ;
      RECT 857.500000 342.350000 858.500000 343.650000 ;
      RECT 816.500000 342.350000 849.500000 343.650000 ;
      RECT 807.500000 342.350000 808.500000 343.650000 ;
      RECT 766.500000 342.350000 799.500000 343.650000 ;
      RECT 757.500000 342.350000 758.500000 343.650000 ;
      RECT 716.500000 342.350000 749.500000 343.650000 ;
      RECT 707.500000 342.350000 708.500000 343.650000 ;
      RECT 666.500000 342.350000 699.500000 343.650000 ;
      RECT 657.500000 342.350000 658.500000 343.650000 ;
      RECT 616.500000 342.350000 649.500000 343.650000 ;
      RECT 607.500000 342.350000 608.500000 343.650000 ;
      RECT 566.500000 342.350000 599.500000 343.650000 ;
      RECT 557.500000 342.350000 558.500000 343.650000 ;
      RECT 516.500000 342.350000 549.500000 343.650000 ;
      RECT 507.500000 342.350000 508.500000 343.650000 ;
      RECT 466.500000 342.350000 499.500000 343.650000 ;
      RECT 457.500000 342.350000 458.500000 343.650000 ;
      RECT 416.500000 342.350000 449.500000 343.650000 ;
      RECT 407.500000 342.350000 408.500000 343.650000 ;
      RECT 366.500000 342.350000 399.500000 343.650000 ;
      RECT 357.500000 342.350000 358.500000 343.650000 ;
      RECT 316.500000 342.350000 349.500000 343.650000 ;
      RECT 307.500000 342.350000 308.500000 343.650000 ;
      RECT 266.500000 342.350000 299.500000 343.650000 ;
      RECT 257.500000 342.350000 258.500000 343.650000 ;
      RECT 216.500000 342.350000 249.500000 343.650000 ;
      RECT 207.500000 342.350000 208.500000 343.650000 ;
      RECT 166.500000 342.350000 199.500000 343.650000 ;
      RECT 157.500000 342.350000 158.500000 343.650000 ;
      RECT 116.500000 342.350000 149.500000 343.650000 ;
      RECT 107.500000 342.350000 108.500000 343.650000 ;
      RECT 66.500000 342.350000 99.500000 343.650000 ;
      RECT 57.500000 342.350000 58.500000 343.650000 ;
      RECT 29.500000 342.350000 49.500000 343.650000 ;
      RECT 15.500000 342.350000 16.500000 343.650000 ;
      RECT 1157.500000 341.650000 1170.500000 342.350000 ;
      RECT 1107.500000 341.650000 1149.500000 342.350000 ;
      RECT 1057.500000 341.650000 1099.500000 342.350000 ;
      RECT 1007.500000 341.650000 1049.500000 342.350000 ;
      RECT 957.500000 341.650000 999.500000 342.350000 ;
      RECT 907.500000 341.650000 949.500000 342.350000 ;
      RECT 857.500000 341.650000 899.500000 342.350000 ;
      RECT 807.500000 341.650000 849.500000 342.350000 ;
      RECT 757.500000 341.650000 799.500000 342.350000 ;
      RECT 707.500000 341.650000 749.500000 342.350000 ;
      RECT 657.500000 341.650000 699.500000 342.350000 ;
      RECT 607.500000 341.650000 649.500000 342.350000 ;
      RECT 557.500000 341.650000 599.500000 342.350000 ;
      RECT 507.500000 341.650000 549.500000 342.350000 ;
      RECT 457.500000 341.650000 499.500000 342.350000 ;
      RECT 407.500000 341.650000 449.500000 342.350000 ;
      RECT 357.500000 341.650000 399.500000 342.350000 ;
      RECT 307.500000 341.650000 349.500000 342.350000 ;
      RECT 257.500000 341.650000 299.500000 342.350000 ;
      RECT 207.500000 341.650000 249.500000 342.350000 ;
      RECT 157.500000 341.650000 199.500000 342.350000 ;
      RECT 107.500000 341.650000 149.500000 342.350000 ;
      RECT 57.500000 341.650000 99.500000 342.350000 ;
      RECT 15.500000 341.650000 49.500000 342.350000 ;
      RECT 1183.500000 340.350000 1186.000000 343.650000 ;
      RECT 1169.500000 340.350000 1170.500000 341.650000 ;
      RECT 1116.500000 340.350000 1149.500000 341.650000 ;
      RECT 1107.500000 340.350000 1108.500000 341.650000 ;
      RECT 1066.500000 340.350000 1099.500000 341.650000 ;
      RECT 1057.500000 340.350000 1058.500000 341.650000 ;
      RECT 1016.500000 340.350000 1049.500000 341.650000 ;
      RECT 1007.500000 340.350000 1008.500000 341.650000 ;
      RECT 966.500000 340.350000 999.500000 341.650000 ;
      RECT 957.500000 340.350000 958.500000 341.650000 ;
      RECT 916.500000 340.350000 949.500000 341.650000 ;
      RECT 907.500000 340.350000 908.500000 341.650000 ;
      RECT 866.500000 340.350000 899.500000 341.650000 ;
      RECT 857.500000 340.350000 858.500000 341.650000 ;
      RECT 816.500000 340.350000 849.500000 341.650000 ;
      RECT 807.500000 340.350000 808.500000 341.650000 ;
      RECT 766.500000 340.350000 799.500000 341.650000 ;
      RECT 757.500000 340.350000 758.500000 341.650000 ;
      RECT 716.500000 340.350000 749.500000 341.650000 ;
      RECT 707.500000 340.350000 708.500000 341.650000 ;
      RECT 666.500000 340.350000 699.500000 341.650000 ;
      RECT 657.500000 340.350000 658.500000 341.650000 ;
      RECT 616.500000 340.350000 649.500000 341.650000 ;
      RECT 607.500000 340.350000 608.500000 341.650000 ;
      RECT 566.500000 340.350000 599.500000 341.650000 ;
      RECT 557.500000 340.350000 558.500000 341.650000 ;
      RECT 516.500000 340.350000 549.500000 341.650000 ;
      RECT 507.500000 340.350000 508.500000 341.650000 ;
      RECT 466.500000 340.350000 499.500000 341.650000 ;
      RECT 457.500000 340.350000 458.500000 341.650000 ;
      RECT 416.500000 340.350000 449.500000 341.650000 ;
      RECT 407.500000 340.350000 408.500000 341.650000 ;
      RECT 366.500000 340.350000 399.500000 341.650000 ;
      RECT 357.500000 340.350000 358.500000 341.650000 ;
      RECT 316.500000 340.350000 349.500000 341.650000 ;
      RECT 307.500000 340.350000 308.500000 341.650000 ;
      RECT 266.500000 340.350000 299.500000 341.650000 ;
      RECT 257.500000 340.350000 258.500000 341.650000 ;
      RECT 216.500000 340.350000 249.500000 341.650000 ;
      RECT 207.500000 340.350000 208.500000 341.650000 ;
      RECT 166.500000 340.350000 199.500000 341.650000 ;
      RECT 157.500000 340.350000 158.500000 341.650000 ;
      RECT 116.500000 340.350000 149.500000 341.650000 ;
      RECT 107.500000 340.350000 108.500000 341.650000 ;
      RECT 66.500000 340.350000 99.500000 341.650000 ;
      RECT 57.500000 340.350000 58.500000 341.650000 ;
      RECT 29.500000 340.350000 49.500000 341.650000 ;
      RECT 15.500000 340.350000 16.500000 341.650000 ;
      RECT 0.000000 340.350000 2.500000 343.650000 ;
      RECT 1169.500000 339.650000 1186.000000 340.350000 ;
      RECT 1116.500000 339.650000 1156.500000 340.350000 ;
      RECT 1066.500000 339.650000 1108.500000 340.350000 ;
      RECT 1016.500000 339.650000 1058.500000 340.350000 ;
      RECT 966.500000 339.650000 1008.500000 340.350000 ;
      RECT 916.500000 339.650000 958.500000 340.350000 ;
      RECT 866.500000 339.650000 908.500000 340.350000 ;
      RECT 816.500000 339.650000 858.500000 340.350000 ;
      RECT 766.500000 339.650000 808.500000 340.350000 ;
      RECT 716.500000 339.650000 758.500000 340.350000 ;
      RECT 666.500000 339.650000 708.500000 340.350000 ;
      RECT 616.500000 339.650000 658.500000 340.350000 ;
      RECT 566.500000 339.650000 608.500000 340.350000 ;
      RECT 516.500000 339.650000 558.500000 340.350000 ;
      RECT 466.500000 339.650000 508.500000 340.350000 ;
      RECT 416.500000 339.650000 458.500000 340.350000 ;
      RECT 366.500000 339.650000 408.500000 340.350000 ;
      RECT 316.500000 339.650000 358.500000 340.350000 ;
      RECT 266.500000 339.650000 308.500000 340.350000 ;
      RECT 216.500000 339.650000 258.500000 340.350000 ;
      RECT 166.500000 339.650000 208.500000 340.350000 ;
      RECT 116.500000 339.650000 158.500000 340.350000 ;
      RECT 66.500000 339.650000 108.500000 340.350000 ;
      RECT 29.500000 339.650000 58.500000 340.350000 ;
      RECT 0.000000 339.650000 16.500000 340.350000 ;
      RECT 1169.500000 338.350000 1170.500000 339.650000 ;
      RECT 1116.500000 338.350000 1149.500000 339.650000 ;
      RECT 1107.500000 338.350000 1108.500000 339.650000 ;
      RECT 1066.500000 338.350000 1099.500000 339.650000 ;
      RECT 1057.500000 338.350000 1058.500000 339.650000 ;
      RECT 1016.500000 338.350000 1049.500000 339.650000 ;
      RECT 1007.500000 338.350000 1008.500000 339.650000 ;
      RECT 966.500000 338.350000 999.500000 339.650000 ;
      RECT 957.500000 338.350000 958.500000 339.650000 ;
      RECT 916.500000 338.350000 949.500000 339.650000 ;
      RECT 907.500000 338.350000 908.500000 339.650000 ;
      RECT 866.500000 338.350000 899.500000 339.650000 ;
      RECT 857.500000 338.350000 858.500000 339.650000 ;
      RECT 816.500000 338.350000 849.500000 339.650000 ;
      RECT 807.500000 338.350000 808.500000 339.650000 ;
      RECT 766.500000 338.350000 799.500000 339.650000 ;
      RECT 757.500000 338.350000 758.500000 339.650000 ;
      RECT 716.500000 338.350000 749.500000 339.650000 ;
      RECT 707.500000 338.350000 708.500000 339.650000 ;
      RECT 666.500000 338.350000 699.500000 339.650000 ;
      RECT 657.500000 338.350000 658.500000 339.650000 ;
      RECT 616.500000 338.350000 649.500000 339.650000 ;
      RECT 607.500000 338.350000 608.500000 339.650000 ;
      RECT 566.500000 338.350000 599.500000 339.650000 ;
      RECT 557.500000 338.350000 558.500000 339.650000 ;
      RECT 516.500000 338.350000 549.500000 339.650000 ;
      RECT 507.500000 338.350000 508.500000 339.650000 ;
      RECT 466.500000 338.350000 499.500000 339.650000 ;
      RECT 457.500000 338.350000 458.500000 339.650000 ;
      RECT 416.500000 338.350000 449.500000 339.650000 ;
      RECT 407.500000 338.350000 408.500000 339.650000 ;
      RECT 366.500000 338.350000 399.500000 339.650000 ;
      RECT 357.500000 338.350000 358.500000 339.650000 ;
      RECT 316.500000 338.350000 349.500000 339.650000 ;
      RECT 307.500000 338.350000 308.500000 339.650000 ;
      RECT 266.500000 338.350000 299.500000 339.650000 ;
      RECT 257.500000 338.350000 258.500000 339.650000 ;
      RECT 216.500000 338.350000 249.500000 339.650000 ;
      RECT 207.500000 338.350000 208.500000 339.650000 ;
      RECT 166.500000 338.350000 199.500000 339.650000 ;
      RECT 157.500000 338.350000 158.500000 339.650000 ;
      RECT 116.500000 338.350000 149.500000 339.650000 ;
      RECT 107.500000 338.350000 108.500000 339.650000 ;
      RECT 66.500000 338.350000 99.500000 339.650000 ;
      RECT 57.500000 338.350000 58.500000 339.650000 ;
      RECT 29.500000 338.350000 49.500000 339.650000 ;
      RECT 15.500000 338.350000 16.500000 339.650000 ;
      RECT 1157.500000 337.650000 1170.500000 338.350000 ;
      RECT 1107.500000 337.650000 1149.500000 338.350000 ;
      RECT 1057.500000 337.650000 1099.500000 338.350000 ;
      RECT 1007.500000 337.650000 1049.500000 338.350000 ;
      RECT 957.500000 337.650000 999.500000 338.350000 ;
      RECT 907.500000 337.650000 949.500000 338.350000 ;
      RECT 857.500000 337.650000 899.500000 338.350000 ;
      RECT 807.500000 337.650000 849.500000 338.350000 ;
      RECT 757.500000 337.650000 799.500000 338.350000 ;
      RECT 707.500000 337.650000 749.500000 338.350000 ;
      RECT 657.500000 337.650000 699.500000 338.350000 ;
      RECT 607.500000 337.650000 649.500000 338.350000 ;
      RECT 557.500000 337.650000 599.500000 338.350000 ;
      RECT 507.500000 337.650000 549.500000 338.350000 ;
      RECT 457.500000 337.650000 499.500000 338.350000 ;
      RECT 407.500000 337.650000 449.500000 338.350000 ;
      RECT 357.500000 337.650000 399.500000 338.350000 ;
      RECT 307.500000 337.650000 349.500000 338.350000 ;
      RECT 257.500000 337.650000 299.500000 338.350000 ;
      RECT 207.500000 337.650000 249.500000 338.350000 ;
      RECT 157.500000 337.650000 199.500000 338.350000 ;
      RECT 107.500000 337.650000 149.500000 338.350000 ;
      RECT 57.500000 337.650000 99.500000 338.350000 ;
      RECT 15.500000 337.650000 49.500000 338.350000 ;
      RECT 1183.500000 336.350000 1186.000000 339.650000 ;
      RECT 1169.500000 336.350000 1170.500000 337.650000 ;
      RECT 1116.500000 336.350000 1149.500000 337.650000 ;
      RECT 1107.500000 336.350000 1108.500000 337.650000 ;
      RECT 1066.500000 336.350000 1099.500000 337.650000 ;
      RECT 1057.500000 336.350000 1058.500000 337.650000 ;
      RECT 1016.500000 336.350000 1049.500000 337.650000 ;
      RECT 1007.500000 336.350000 1008.500000 337.650000 ;
      RECT 966.500000 336.350000 999.500000 337.650000 ;
      RECT 957.500000 336.350000 958.500000 337.650000 ;
      RECT 916.500000 336.350000 949.500000 337.650000 ;
      RECT 907.500000 336.350000 908.500000 337.650000 ;
      RECT 866.500000 336.350000 899.500000 337.650000 ;
      RECT 857.500000 336.350000 858.500000 337.650000 ;
      RECT 816.500000 336.350000 849.500000 337.650000 ;
      RECT 807.500000 336.350000 808.500000 337.650000 ;
      RECT 766.500000 336.350000 799.500000 337.650000 ;
      RECT 757.500000 336.350000 758.500000 337.650000 ;
      RECT 716.500000 336.350000 749.500000 337.650000 ;
      RECT 707.500000 336.350000 708.500000 337.650000 ;
      RECT 666.500000 336.350000 699.500000 337.650000 ;
      RECT 657.500000 336.350000 658.500000 337.650000 ;
      RECT 616.500000 336.350000 649.500000 337.650000 ;
      RECT 607.500000 336.350000 608.500000 337.650000 ;
      RECT 566.500000 336.350000 599.500000 337.650000 ;
      RECT 557.500000 336.350000 558.500000 337.650000 ;
      RECT 516.500000 336.350000 549.500000 337.650000 ;
      RECT 507.500000 336.350000 508.500000 337.650000 ;
      RECT 466.500000 336.350000 499.500000 337.650000 ;
      RECT 457.500000 336.350000 458.500000 337.650000 ;
      RECT 416.500000 336.350000 449.500000 337.650000 ;
      RECT 407.500000 336.350000 408.500000 337.650000 ;
      RECT 366.500000 336.350000 399.500000 337.650000 ;
      RECT 357.500000 336.350000 358.500000 337.650000 ;
      RECT 316.500000 336.350000 349.500000 337.650000 ;
      RECT 307.500000 336.350000 308.500000 337.650000 ;
      RECT 266.500000 336.350000 299.500000 337.650000 ;
      RECT 257.500000 336.350000 258.500000 337.650000 ;
      RECT 216.500000 336.350000 249.500000 337.650000 ;
      RECT 207.500000 336.350000 208.500000 337.650000 ;
      RECT 166.500000 336.350000 199.500000 337.650000 ;
      RECT 157.500000 336.350000 158.500000 337.650000 ;
      RECT 116.500000 336.350000 149.500000 337.650000 ;
      RECT 107.500000 336.350000 108.500000 337.650000 ;
      RECT 66.500000 336.350000 99.500000 337.650000 ;
      RECT 57.500000 336.350000 58.500000 337.650000 ;
      RECT 29.500000 336.350000 49.500000 337.650000 ;
      RECT 15.500000 336.350000 16.500000 337.650000 ;
      RECT 0.000000 336.350000 2.500000 339.650000 ;
      RECT 1169.500000 335.650000 1186.000000 336.350000 ;
      RECT 1116.500000 335.650000 1156.500000 336.350000 ;
      RECT 1066.500000 335.650000 1108.500000 336.350000 ;
      RECT 1016.500000 335.650000 1058.500000 336.350000 ;
      RECT 966.500000 335.650000 1008.500000 336.350000 ;
      RECT 916.500000 335.650000 958.500000 336.350000 ;
      RECT 866.500000 335.650000 908.500000 336.350000 ;
      RECT 816.500000 335.650000 858.500000 336.350000 ;
      RECT 766.500000 335.650000 808.500000 336.350000 ;
      RECT 716.500000 335.650000 758.500000 336.350000 ;
      RECT 666.500000 335.650000 708.500000 336.350000 ;
      RECT 616.500000 335.650000 658.500000 336.350000 ;
      RECT 566.500000 335.650000 608.500000 336.350000 ;
      RECT 516.500000 335.650000 558.500000 336.350000 ;
      RECT 466.500000 335.650000 508.500000 336.350000 ;
      RECT 416.500000 335.650000 458.500000 336.350000 ;
      RECT 366.500000 335.650000 408.500000 336.350000 ;
      RECT 316.500000 335.650000 358.500000 336.350000 ;
      RECT 266.500000 335.650000 308.500000 336.350000 ;
      RECT 216.500000 335.650000 258.500000 336.350000 ;
      RECT 166.500000 335.650000 208.500000 336.350000 ;
      RECT 116.500000 335.650000 158.500000 336.350000 ;
      RECT 66.500000 335.650000 108.500000 336.350000 ;
      RECT 29.500000 335.650000 58.500000 336.350000 ;
      RECT 0.000000 335.650000 16.500000 336.350000 ;
      RECT 1169.500000 334.350000 1170.500000 335.650000 ;
      RECT 1116.500000 334.350000 1149.500000 335.650000 ;
      RECT 1107.500000 334.350000 1108.500000 335.650000 ;
      RECT 1066.500000 334.350000 1099.500000 335.650000 ;
      RECT 1057.500000 334.350000 1058.500000 335.650000 ;
      RECT 1016.500000 334.350000 1049.500000 335.650000 ;
      RECT 1007.500000 334.350000 1008.500000 335.650000 ;
      RECT 966.500000 334.350000 999.500000 335.650000 ;
      RECT 957.500000 334.350000 958.500000 335.650000 ;
      RECT 916.500000 334.350000 949.500000 335.650000 ;
      RECT 907.500000 334.350000 908.500000 335.650000 ;
      RECT 866.500000 334.350000 899.500000 335.650000 ;
      RECT 857.500000 334.350000 858.500000 335.650000 ;
      RECT 816.500000 334.350000 849.500000 335.650000 ;
      RECT 807.500000 334.350000 808.500000 335.650000 ;
      RECT 766.500000 334.350000 799.500000 335.650000 ;
      RECT 757.500000 334.350000 758.500000 335.650000 ;
      RECT 716.500000 334.350000 749.500000 335.650000 ;
      RECT 707.500000 334.350000 708.500000 335.650000 ;
      RECT 666.500000 334.350000 699.500000 335.650000 ;
      RECT 657.500000 334.350000 658.500000 335.650000 ;
      RECT 616.500000 334.350000 649.500000 335.650000 ;
      RECT 607.500000 334.350000 608.500000 335.650000 ;
      RECT 566.500000 334.350000 599.500000 335.650000 ;
      RECT 557.500000 334.350000 558.500000 335.650000 ;
      RECT 516.500000 334.350000 549.500000 335.650000 ;
      RECT 507.500000 334.350000 508.500000 335.650000 ;
      RECT 466.500000 334.350000 499.500000 335.650000 ;
      RECT 457.500000 334.350000 458.500000 335.650000 ;
      RECT 416.500000 334.350000 449.500000 335.650000 ;
      RECT 407.500000 334.350000 408.500000 335.650000 ;
      RECT 366.500000 334.350000 399.500000 335.650000 ;
      RECT 357.500000 334.350000 358.500000 335.650000 ;
      RECT 316.500000 334.350000 349.500000 335.650000 ;
      RECT 307.500000 334.350000 308.500000 335.650000 ;
      RECT 266.500000 334.350000 299.500000 335.650000 ;
      RECT 257.500000 334.350000 258.500000 335.650000 ;
      RECT 216.500000 334.350000 249.500000 335.650000 ;
      RECT 207.500000 334.350000 208.500000 335.650000 ;
      RECT 166.500000 334.350000 199.500000 335.650000 ;
      RECT 157.500000 334.350000 158.500000 335.650000 ;
      RECT 116.500000 334.350000 149.500000 335.650000 ;
      RECT 107.500000 334.350000 108.500000 335.650000 ;
      RECT 66.500000 334.350000 99.500000 335.650000 ;
      RECT 57.500000 334.350000 58.500000 335.650000 ;
      RECT 29.500000 334.350000 49.500000 335.650000 ;
      RECT 15.500000 334.350000 16.500000 335.650000 ;
      RECT 1157.500000 333.650000 1170.500000 334.350000 ;
      RECT 1107.500000 333.650000 1149.500000 334.350000 ;
      RECT 1057.500000 333.650000 1099.500000 334.350000 ;
      RECT 1007.500000 333.650000 1049.500000 334.350000 ;
      RECT 957.500000 333.650000 999.500000 334.350000 ;
      RECT 907.500000 333.650000 949.500000 334.350000 ;
      RECT 857.500000 333.650000 899.500000 334.350000 ;
      RECT 807.500000 333.650000 849.500000 334.350000 ;
      RECT 757.500000 333.650000 799.500000 334.350000 ;
      RECT 707.500000 333.650000 749.500000 334.350000 ;
      RECT 657.500000 333.650000 699.500000 334.350000 ;
      RECT 607.500000 333.650000 649.500000 334.350000 ;
      RECT 557.500000 333.650000 599.500000 334.350000 ;
      RECT 507.500000 333.650000 549.500000 334.350000 ;
      RECT 457.500000 333.650000 499.500000 334.350000 ;
      RECT 407.500000 333.650000 449.500000 334.350000 ;
      RECT 357.500000 333.650000 399.500000 334.350000 ;
      RECT 307.500000 333.650000 349.500000 334.350000 ;
      RECT 257.500000 333.650000 299.500000 334.350000 ;
      RECT 207.500000 333.650000 249.500000 334.350000 ;
      RECT 157.500000 333.650000 199.500000 334.350000 ;
      RECT 107.500000 333.650000 149.500000 334.350000 ;
      RECT 57.500000 333.650000 99.500000 334.350000 ;
      RECT 15.500000 333.650000 49.500000 334.350000 ;
      RECT 1183.500000 332.350000 1186.000000 335.650000 ;
      RECT 1169.500000 332.350000 1170.500000 333.650000 ;
      RECT 1116.500000 332.350000 1149.500000 333.650000 ;
      RECT 1107.500000 332.350000 1108.500000 333.650000 ;
      RECT 1066.500000 332.350000 1099.500000 333.650000 ;
      RECT 1057.500000 332.350000 1058.500000 333.650000 ;
      RECT 1016.500000 332.350000 1049.500000 333.650000 ;
      RECT 1007.500000 332.350000 1008.500000 333.650000 ;
      RECT 966.500000 332.350000 999.500000 333.650000 ;
      RECT 957.500000 332.350000 958.500000 333.650000 ;
      RECT 916.500000 332.350000 949.500000 333.650000 ;
      RECT 907.500000 332.350000 908.500000 333.650000 ;
      RECT 866.500000 332.350000 899.500000 333.650000 ;
      RECT 857.500000 332.350000 858.500000 333.650000 ;
      RECT 816.500000 332.350000 849.500000 333.650000 ;
      RECT 807.500000 332.350000 808.500000 333.650000 ;
      RECT 766.500000 332.350000 799.500000 333.650000 ;
      RECT 757.500000 332.350000 758.500000 333.650000 ;
      RECT 716.500000 332.350000 749.500000 333.650000 ;
      RECT 707.500000 332.350000 708.500000 333.650000 ;
      RECT 666.500000 332.350000 699.500000 333.650000 ;
      RECT 657.500000 332.350000 658.500000 333.650000 ;
      RECT 616.500000 332.350000 649.500000 333.650000 ;
      RECT 607.500000 332.350000 608.500000 333.650000 ;
      RECT 566.500000 332.350000 599.500000 333.650000 ;
      RECT 557.500000 332.350000 558.500000 333.650000 ;
      RECT 516.500000 332.350000 549.500000 333.650000 ;
      RECT 507.500000 332.350000 508.500000 333.650000 ;
      RECT 466.500000 332.350000 499.500000 333.650000 ;
      RECT 457.500000 332.350000 458.500000 333.650000 ;
      RECT 416.500000 332.350000 449.500000 333.650000 ;
      RECT 407.500000 332.350000 408.500000 333.650000 ;
      RECT 366.500000 332.350000 399.500000 333.650000 ;
      RECT 357.500000 332.350000 358.500000 333.650000 ;
      RECT 316.500000 332.350000 349.500000 333.650000 ;
      RECT 307.500000 332.350000 308.500000 333.650000 ;
      RECT 266.500000 332.350000 299.500000 333.650000 ;
      RECT 257.500000 332.350000 258.500000 333.650000 ;
      RECT 216.500000 332.350000 249.500000 333.650000 ;
      RECT 207.500000 332.350000 208.500000 333.650000 ;
      RECT 166.500000 332.350000 199.500000 333.650000 ;
      RECT 157.500000 332.350000 158.500000 333.650000 ;
      RECT 116.500000 332.350000 149.500000 333.650000 ;
      RECT 107.500000 332.350000 108.500000 333.650000 ;
      RECT 66.500000 332.350000 99.500000 333.650000 ;
      RECT 57.500000 332.350000 58.500000 333.650000 ;
      RECT 29.500000 332.350000 49.500000 333.650000 ;
      RECT 15.500000 332.350000 16.500000 333.650000 ;
      RECT 0.000000 332.350000 2.500000 335.650000 ;
      RECT 1169.500000 331.650000 1186.000000 332.350000 ;
      RECT 1116.500000 331.650000 1156.500000 332.350000 ;
      RECT 1066.500000 331.650000 1108.500000 332.350000 ;
      RECT 1016.500000 331.650000 1058.500000 332.350000 ;
      RECT 966.500000 331.650000 1008.500000 332.350000 ;
      RECT 916.500000 331.650000 958.500000 332.350000 ;
      RECT 866.500000 331.650000 908.500000 332.350000 ;
      RECT 816.500000 331.650000 858.500000 332.350000 ;
      RECT 766.500000 331.650000 808.500000 332.350000 ;
      RECT 716.500000 331.650000 758.500000 332.350000 ;
      RECT 666.500000 331.650000 708.500000 332.350000 ;
      RECT 616.500000 331.650000 658.500000 332.350000 ;
      RECT 566.500000 331.650000 608.500000 332.350000 ;
      RECT 516.500000 331.650000 558.500000 332.350000 ;
      RECT 466.500000 331.650000 508.500000 332.350000 ;
      RECT 416.500000 331.650000 458.500000 332.350000 ;
      RECT 366.500000 331.650000 408.500000 332.350000 ;
      RECT 316.500000 331.650000 358.500000 332.350000 ;
      RECT 266.500000 331.650000 308.500000 332.350000 ;
      RECT 216.500000 331.650000 258.500000 332.350000 ;
      RECT 166.500000 331.650000 208.500000 332.350000 ;
      RECT 116.500000 331.650000 158.500000 332.350000 ;
      RECT 66.500000 331.650000 108.500000 332.350000 ;
      RECT 29.500000 331.650000 58.500000 332.350000 ;
      RECT 0.000000 331.650000 16.500000 332.350000 ;
      RECT 1169.500000 330.350000 1170.500000 331.650000 ;
      RECT 1116.500000 330.350000 1149.500000 331.650000 ;
      RECT 1107.500000 330.350000 1108.500000 331.650000 ;
      RECT 1066.500000 330.350000 1099.500000 331.650000 ;
      RECT 1057.500000 330.350000 1058.500000 331.650000 ;
      RECT 1016.500000 330.350000 1049.500000 331.650000 ;
      RECT 1007.500000 330.350000 1008.500000 331.650000 ;
      RECT 966.500000 330.350000 999.500000 331.650000 ;
      RECT 957.500000 330.350000 958.500000 331.650000 ;
      RECT 916.500000 330.350000 949.500000 331.650000 ;
      RECT 907.500000 330.350000 908.500000 331.650000 ;
      RECT 866.500000 330.350000 899.500000 331.650000 ;
      RECT 857.500000 330.350000 858.500000 331.650000 ;
      RECT 816.500000 330.350000 849.500000 331.650000 ;
      RECT 807.500000 330.350000 808.500000 331.650000 ;
      RECT 766.500000 330.350000 799.500000 331.650000 ;
      RECT 757.500000 330.350000 758.500000 331.650000 ;
      RECT 716.500000 330.350000 749.500000 331.650000 ;
      RECT 707.500000 330.350000 708.500000 331.650000 ;
      RECT 666.500000 330.350000 699.500000 331.650000 ;
      RECT 657.500000 330.350000 658.500000 331.650000 ;
      RECT 616.500000 330.350000 649.500000 331.650000 ;
      RECT 607.500000 330.350000 608.500000 331.650000 ;
      RECT 566.500000 330.350000 599.500000 331.650000 ;
      RECT 557.500000 330.350000 558.500000 331.650000 ;
      RECT 516.500000 330.350000 549.500000 331.650000 ;
      RECT 507.500000 330.350000 508.500000 331.650000 ;
      RECT 466.500000 330.350000 499.500000 331.650000 ;
      RECT 457.500000 330.350000 458.500000 331.650000 ;
      RECT 416.500000 330.350000 449.500000 331.650000 ;
      RECT 407.500000 330.350000 408.500000 331.650000 ;
      RECT 366.500000 330.350000 399.500000 331.650000 ;
      RECT 357.500000 330.350000 358.500000 331.650000 ;
      RECT 316.500000 330.350000 349.500000 331.650000 ;
      RECT 307.500000 330.350000 308.500000 331.650000 ;
      RECT 266.500000 330.350000 299.500000 331.650000 ;
      RECT 257.500000 330.350000 258.500000 331.650000 ;
      RECT 216.500000 330.350000 249.500000 331.650000 ;
      RECT 207.500000 330.350000 208.500000 331.650000 ;
      RECT 166.500000 330.350000 199.500000 331.650000 ;
      RECT 157.500000 330.350000 158.500000 331.650000 ;
      RECT 116.500000 330.350000 149.500000 331.650000 ;
      RECT 107.500000 330.350000 108.500000 331.650000 ;
      RECT 66.500000 330.350000 99.500000 331.650000 ;
      RECT 57.500000 330.350000 58.500000 331.650000 ;
      RECT 29.500000 330.350000 49.500000 331.650000 ;
      RECT 15.500000 330.350000 16.500000 331.650000 ;
      RECT 1157.500000 329.650000 1170.500000 330.350000 ;
      RECT 1107.500000 329.650000 1149.500000 330.350000 ;
      RECT 1057.500000 329.650000 1099.500000 330.350000 ;
      RECT 1007.500000 329.650000 1049.500000 330.350000 ;
      RECT 957.500000 329.650000 999.500000 330.350000 ;
      RECT 907.500000 329.650000 949.500000 330.350000 ;
      RECT 857.500000 329.650000 899.500000 330.350000 ;
      RECT 807.500000 329.650000 849.500000 330.350000 ;
      RECT 757.500000 329.650000 799.500000 330.350000 ;
      RECT 707.500000 329.650000 749.500000 330.350000 ;
      RECT 657.500000 329.650000 699.500000 330.350000 ;
      RECT 607.500000 329.650000 649.500000 330.350000 ;
      RECT 557.500000 329.650000 599.500000 330.350000 ;
      RECT 507.500000 329.650000 549.500000 330.350000 ;
      RECT 457.500000 329.650000 499.500000 330.350000 ;
      RECT 407.500000 329.650000 449.500000 330.350000 ;
      RECT 357.500000 329.650000 399.500000 330.350000 ;
      RECT 307.500000 329.650000 349.500000 330.350000 ;
      RECT 257.500000 329.650000 299.500000 330.350000 ;
      RECT 207.500000 329.650000 249.500000 330.350000 ;
      RECT 157.500000 329.650000 199.500000 330.350000 ;
      RECT 107.500000 329.650000 149.500000 330.350000 ;
      RECT 57.500000 329.650000 99.500000 330.350000 ;
      RECT 15.500000 329.650000 49.500000 330.350000 ;
      RECT 1183.500000 328.350000 1186.000000 331.650000 ;
      RECT 1169.500000 328.350000 1170.500000 329.650000 ;
      RECT 1116.500000 328.350000 1149.500000 329.650000 ;
      RECT 1107.500000 328.350000 1108.500000 329.650000 ;
      RECT 1066.500000 328.350000 1099.500000 329.650000 ;
      RECT 1057.500000 328.350000 1058.500000 329.650000 ;
      RECT 1016.500000 328.350000 1049.500000 329.650000 ;
      RECT 1007.500000 328.350000 1008.500000 329.650000 ;
      RECT 966.500000 328.350000 999.500000 329.650000 ;
      RECT 957.500000 328.350000 958.500000 329.650000 ;
      RECT 916.500000 328.350000 949.500000 329.650000 ;
      RECT 907.500000 328.350000 908.500000 329.650000 ;
      RECT 866.500000 328.350000 899.500000 329.650000 ;
      RECT 857.500000 328.350000 858.500000 329.650000 ;
      RECT 816.500000 328.350000 849.500000 329.650000 ;
      RECT 807.500000 328.350000 808.500000 329.650000 ;
      RECT 766.500000 328.350000 799.500000 329.650000 ;
      RECT 757.500000 328.350000 758.500000 329.650000 ;
      RECT 716.500000 328.350000 749.500000 329.650000 ;
      RECT 707.500000 328.350000 708.500000 329.650000 ;
      RECT 666.500000 328.350000 699.500000 329.650000 ;
      RECT 657.500000 328.350000 658.500000 329.650000 ;
      RECT 616.500000 328.350000 649.500000 329.650000 ;
      RECT 607.500000 328.350000 608.500000 329.650000 ;
      RECT 566.500000 328.350000 599.500000 329.650000 ;
      RECT 557.500000 328.350000 558.500000 329.650000 ;
      RECT 516.500000 328.350000 549.500000 329.650000 ;
      RECT 507.500000 328.350000 508.500000 329.650000 ;
      RECT 466.500000 328.350000 499.500000 329.650000 ;
      RECT 457.500000 328.350000 458.500000 329.650000 ;
      RECT 416.500000 328.350000 449.500000 329.650000 ;
      RECT 407.500000 328.350000 408.500000 329.650000 ;
      RECT 366.500000 328.350000 399.500000 329.650000 ;
      RECT 357.500000 328.350000 358.500000 329.650000 ;
      RECT 316.500000 328.350000 349.500000 329.650000 ;
      RECT 307.500000 328.350000 308.500000 329.650000 ;
      RECT 266.500000 328.350000 299.500000 329.650000 ;
      RECT 257.500000 328.350000 258.500000 329.650000 ;
      RECT 216.500000 328.350000 249.500000 329.650000 ;
      RECT 207.500000 328.350000 208.500000 329.650000 ;
      RECT 166.500000 328.350000 199.500000 329.650000 ;
      RECT 157.500000 328.350000 158.500000 329.650000 ;
      RECT 116.500000 328.350000 149.500000 329.650000 ;
      RECT 107.500000 328.350000 108.500000 329.650000 ;
      RECT 66.500000 328.350000 99.500000 329.650000 ;
      RECT 57.500000 328.350000 58.500000 329.650000 ;
      RECT 29.500000 328.350000 49.500000 329.650000 ;
      RECT 15.500000 328.350000 16.500000 329.650000 ;
      RECT 0.000000 328.350000 2.500000 331.650000 ;
      RECT 1169.500000 327.650000 1186.000000 328.350000 ;
      RECT 1116.500000 327.650000 1156.500000 328.350000 ;
      RECT 1066.500000 327.650000 1108.500000 328.350000 ;
      RECT 1016.500000 327.650000 1058.500000 328.350000 ;
      RECT 966.500000 327.650000 1008.500000 328.350000 ;
      RECT 916.500000 327.650000 958.500000 328.350000 ;
      RECT 866.500000 327.650000 908.500000 328.350000 ;
      RECT 816.500000 327.650000 858.500000 328.350000 ;
      RECT 766.500000 327.650000 808.500000 328.350000 ;
      RECT 716.500000 327.650000 758.500000 328.350000 ;
      RECT 666.500000 327.650000 708.500000 328.350000 ;
      RECT 616.500000 327.650000 658.500000 328.350000 ;
      RECT 566.500000 327.650000 608.500000 328.350000 ;
      RECT 516.500000 327.650000 558.500000 328.350000 ;
      RECT 466.500000 327.650000 508.500000 328.350000 ;
      RECT 416.500000 327.650000 458.500000 328.350000 ;
      RECT 366.500000 327.650000 408.500000 328.350000 ;
      RECT 316.500000 327.650000 358.500000 328.350000 ;
      RECT 266.500000 327.650000 308.500000 328.350000 ;
      RECT 216.500000 327.650000 258.500000 328.350000 ;
      RECT 166.500000 327.650000 208.500000 328.350000 ;
      RECT 116.500000 327.650000 158.500000 328.350000 ;
      RECT 66.500000 327.650000 108.500000 328.350000 ;
      RECT 29.500000 327.650000 58.500000 328.350000 ;
      RECT 0.000000 327.650000 16.500000 328.350000 ;
      RECT 1169.500000 326.350000 1170.500000 327.650000 ;
      RECT 1116.500000 326.350000 1149.500000 327.650000 ;
      RECT 1107.500000 326.350000 1108.500000 327.650000 ;
      RECT 1066.500000 326.350000 1099.500000 327.650000 ;
      RECT 1057.500000 326.350000 1058.500000 327.650000 ;
      RECT 1016.500000 326.350000 1049.500000 327.650000 ;
      RECT 1007.500000 326.350000 1008.500000 327.650000 ;
      RECT 966.500000 326.350000 999.500000 327.650000 ;
      RECT 957.500000 326.350000 958.500000 327.650000 ;
      RECT 916.500000 326.350000 949.500000 327.650000 ;
      RECT 907.500000 326.350000 908.500000 327.650000 ;
      RECT 866.500000 326.350000 899.500000 327.650000 ;
      RECT 857.500000 326.350000 858.500000 327.650000 ;
      RECT 816.500000 326.350000 849.500000 327.650000 ;
      RECT 807.500000 326.350000 808.500000 327.650000 ;
      RECT 766.500000 326.350000 799.500000 327.650000 ;
      RECT 757.500000 326.350000 758.500000 327.650000 ;
      RECT 716.500000 326.350000 749.500000 327.650000 ;
      RECT 707.500000 326.350000 708.500000 327.650000 ;
      RECT 666.500000 326.350000 699.500000 327.650000 ;
      RECT 657.500000 326.350000 658.500000 327.650000 ;
      RECT 616.500000 326.350000 649.500000 327.650000 ;
      RECT 607.500000 326.350000 608.500000 327.650000 ;
      RECT 566.500000 326.350000 599.500000 327.650000 ;
      RECT 557.500000 326.350000 558.500000 327.650000 ;
      RECT 516.500000 326.350000 549.500000 327.650000 ;
      RECT 507.500000 326.350000 508.500000 327.650000 ;
      RECT 466.500000 326.350000 499.500000 327.650000 ;
      RECT 457.500000 326.350000 458.500000 327.650000 ;
      RECT 416.500000 326.350000 449.500000 327.650000 ;
      RECT 407.500000 326.350000 408.500000 327.650000 ;
      RECT 366.500000 326.350000 399.500000 327.650000 ;
      RECT 357.500000 326.350000 358.500000 327.650000 ;
      RECT 316.500000 326.350000 349.500000 327.650000 ;
      RECT 307.500000 326.350000 308.500000 327.650000 ;
      RECT 266.500000 326.350000 299.500000 327.650000 ;
      RECT 257.500000 326.350000 258.500000 327.650000 ;
      RECT 216.500000 326.350000 249.500000 327.650000 ;
      RECT 207.500000 326.350000 208.500000 327.650000 ;
      RECT 166.500000 326.350000 199.500000 327.650000 ;
      RECT 157.500000 326.350000 158.500000 327.650000 ;
      RECT 116.500000 326.350000 149.500000 327.650000 ;
      RECT 107.500000 326.350000 108.500000 327.650000 ;
      RECT 66.500000 326.350000 99.500000 327.650000 ;
      RECT 57.500000 326.350000 58.500000 327.650000 ;
      RECT 29.500000 326.350000 49.500000 327.650000 ;
      RECT 15.500000 326.350000 16.500000 327.650000 ;
      RECT 1157.500000 325.650000 1170.500000 326.350000 ;
      RECT 1107.500000 325.650000 1149.500000 326.350000 ;
      RECT 1057.500000 325.650000 1099.500000 326.350000 ;
      RECT 1007.500000 325.650000 1049.500000 326.350000 ;
      RECT 957.500000 325.650000 999.500000 326.350000 ;
      RECT 907.500000 325.650000 949.500000 326.350000 ;
      RECT 857.500000 325.650000 899.500000 326.350000 ;
      RECT 807.500000 325.650000 849.500000 326.350000 ;
      RECT 757.500000 325.650000 799.500000 326.350000 ;
      RECT 707.500000 325.650000 749.500000 326.350000 ;
      RECT 657.500000 325.650000 699.500000 326.350000 ;
      RECT 607.500000 325.650000 649.500000 326.350000 ;
      RECT 557.500000 325.650000 599.500000 326.350000 ;
      RECT 507.500000 325.650000 549.500000 326.350000 ;
      RECT 457.500000 325.650000 499.500000 326.350000 ;
      RECT 407.500000 325.650000 449.500000 326.350000 ;
      RECT 357.500000 325.650000 399.500000 326.350000 ;
      RECT 307.500000 325.650000 349.500000 326.350000 ;
      RECT 257.500000 325.650000 299.500000 326.350000 ;
      RECT 207.500000 325.650000 249.500000 326.350000 ;
      RECT 157.500000 325.650000 199.500000 326.350000 ;
      RECT 107.500000 325.650000 149.500000 326.350000 ;
      RECT 57.500000 325.650000 99.500000 326.350000 ;
      RECT 15.500000 325.650000 49.500000 326.350000 ;
      RECT 1183.500000 324.350000 1186.000000 327.650000 ;
      RECT 1169.500000 324.350000 1170.500000 325.650000 ;
      RECT 1116.500000 324.350000 1149.500000 325.650000 ;
      RECT 1107.500000 324.350000 1108.500000 325.650000 ;
      RECT 1066.500000 324.350000 1099.500000 325.650000 ;
      RECT 1057.500000 324.350000 1058.500000 325.650000 ;
      RECT 1016.500000 324.350000 1049.500000 325.650000 ;
      RECT 1007.500000 324.350000 1008.500000 325.650000 ;
      RECT 966.500000 324.350000 999.500000 325.650000 ;
      RECT 957.500000 324.350000 958.500000 325.650000 ;
      RECT 916.500000 324.350000 949.500000 325.650000 ;
      RECT 907.500000 324.350000 908.500000 325.650000 ;
      RECT 866.500000 324.350000 899.500000 325.650000 ;
      RECT 857.500000 324.350000 858.500000 325.650000 ;
      RECT 816.500000 324.350000 849.500000 325.650000 ;
      RECT 807.500000 324.350000 808.500000 325.650000 ;
      RECT 766.500000 324.350000 799.500000 325.650000 ;
      RECT 757.500000 324.350000 758.500000 325.650000 ;
      RECT 716.500000 324.350000 749.500000 325.650000 ;
      RECT 707.500000 324.350000 708.500000 325.650000 ;
      RECT 666.500000 324.350000 699.500000 325.650000 ;
      RECT 657.500000 324.350000 658.500000 325.650000 ;
      RECT 616.500000 324.350000 649.500000 325.650000 ;
      RECT 607.500000 324.350000 608.500000 325.650000 ;
      RECT 566.500000 324.350000 599.500000 325.650000 ;
      RECT 557.500000 324.350000 558.500000 325.650000 ;
      RECT 516.500000 324.350000 549.500000 325.650000 ;
      RECT 507.500000 324.350000 508.500000 325.650000 ;
      RECT 466.500000 324.350000 499.500000 325.650000 ;
      RECT 457.500000 324.350000 458.500000 325.650000 ;
      RECT 416.500000 324.350000 449.500000 325.650000 ;
      RECT 407.500000 324.350000 408.500000 325.650000 ;
      RECT 366.500000 324.350000 399.500000 325.650000 ;
      RECT 357.500000 324.350000 358.500000 325.650000 ;
      RECT 316.500000 324.350000 349.500000 325.650000 ;
      RECT 307.500000 324.350000 308.500000 325.650000 ;
      RECT 266.500000 324.350000 299.500000 325.650000 ;
      RECT 257.500000 324.350000 258.500000 325.650000 ;
      RECT 216.500000 324.350000 249.500000 325.650000 ;
      RECT 207.500000 324.350000 208.500000 325.650000 ;
      RECT 166.500000 324.350000 199.500000 325.650000 ;
      RECT 157.500000 324.350000 158.500000 325.650000 ;
      RECT 116.500000 324.350000 149.500000 325.650000 ;
      RECT 107.500000 324.350000 108.500000 325.650000 ;
      RECT 66.500000 324.350000 99.500000 325.650000 ;
      RECT 57.500000 324.350000 58.500000 325.650000 ;
      RECT 29.500000 324.350000 49.500000 325.650000 ;
      RECT 15.500000 324.350000 16.500000 325.650000 ;
      RECT 0.000000 324.350000 2.500000 327.650000 ;
      RECT 1169.500000 323.650000 1186.000000 324.350000 ;
      RECT 1116.500000 323.650000 1156.500000 324.350000 ;
      RECT 1066.500000 323.650000 1108.500000 324.350000 ;
      RECT 1016.500000 323.650000 1058.500000 324.350000 ;
      RECT 966.500000 323.650000 1008.500000 324.350000 ;
      RECT 916.500000 323.650000 958.500000 324.350000 ;
      RECT 866.500000 323.650000 908.500000 324.350000 ;
      RECT 816.500000 323.650000 858.500000 324.350000 ;
      RECT 766.500000 323.650000 808.500000 324.350000 ;
      RECT 716.500000 323.650000 758.500000 324.350000 ;
      RECT 666.500000 323.650000 708.500000 324.350000 ;
      RECT 616.500000 323.650000 658.500000 324.350000 ;
      RECT 566.500000 323.650000 608.500000 324.350000 ;
      RECT 516.500000 323.650000 558.500000 324.350000 ;
      RECT 466.500000 323.650000 508.500000 324.350000 ;
      RECT 416.500000 323.650000 458.500000 324.350000 ;
      RECT 366.500000 323.650000 408.500000 324.350000 ;
      RECT 316.500000 323.650000 358.500000 324.350000 ;
      RECT 266.500000 323.650000 308.500000 324.350000 ;
      RECT 216.500000 323.650000 258.500000 324.350000 ;
      RECT 166.500000 323.650000 208.500000 324.350000 ;
      RECT 116.500000 323.650000 158.500000 324.350000 ;
      RECT 66.500000 323.650000 108.500000 324.350000 ;
      RECT 29.500000 323.650000 58.500000 324.350000 ;
      RECT 0.000000 323.650000 16.500000 324.350000 ;
      RECT 1169.500000 322.350000 1170.500000 323.650000 ;
      RECT 1116.500000 322.350000 1149.500000 323.650000 ;
      RECT 1107.500000 322.350000 1108.500000 323.650000 ;
      RECT 1066.500000 322.350000 1099.500000 323.650000 ;
      RECT 1057.500000 322.350000 1058.500000 323.650000 ;
      RECT 1016.500000 322.350000 1049.500000 323.650000 ;
      RECT 1007.500000 322.350000 1008.500000 323.650000 ;
      RECT 966.500000 322.350000 999.500000 323.650000 ;
      RECT 957.500000 322.350000 958.500000 323.650000 ;
      RECT 916.500000 322.350000 949.500000 323.650000 ;
      RECT 907.500000 322.350000 908.500000 323.650000 ;
      RECT 866.500000 322.350000 899.500000 323.650000 ;
      RECT 857.500000 322.350000 858.500000 323.650000 ;
      RECT 816.500000 322.350000 849.500000 323.650000 ;
      RECT 807.500000 322.350000 808.500000 323.650000 ;
      RECT 766.500000 322.350000 799.500000 323.650000 ;
      RECT 757.500000 322.350000 758.500000 323.650000 ;
      RECT 716.500000 322.350000 749.500000 323.650000 ;
      RECT 707.500000 322.350000 708.500000 323.650000 ;
      RECT 666.500000 322.350000 699.500000 323.650000 ;
      RECT 657.500000 322.350000 658.500000 323.650000 ;
      RECT 616.500000 322.350000 649.500000 323.650000 ;
      RECT 607.500000 322.350000 608.500000 323.650000 ;
      RECT 566.500000 322.350000 599.500000 323.650000 ;
      RECT 557.500000 322.350000 558.500000 323.650000 ;
      RECT 516.500000 322.350000 549.500000 323.650000 ;
      RECT 507.500000 322.350000 508.500000 323.650000 ;
      RECT 466.500000 322.350000 499.500000 323.650000 ;
      RECT 457.500000 322.350000 458.500000 323.650000 ;
      RECT 416.500000 322.350000 449.500000 323.650000 ;
      RECT 407.500000 322.350000 408.500000 323.650000 ;
      RECT 366.500000 322.350000 399.500000 323.650000 ;
      RECT 357.500000 322.350000 358.500000 323.650000 ;
      RECT 316.500000 322.350000 349.500000 323.650000 ;
      RECT 307.500000 322.350000 308.500000 323.650000 ;
      RECT 266.500000 322.350000 299.500000 323.650000 ;
      RECT 257.500000 322.350000 258.500000 323.650000 ;
      RECT 216.500000 322.350000 249.500000 323.650000 ;
      RECT 207.500000 322.350000 208.500000 323.650000 ;
      RECT 166.500000 322.350000 199.500000 323.650000 ;
      RECT 157.500000 322.350000 158.500000 323.650000 ;
      RECT 116.500000 322.350000 149.500000 323.650000 ;
      RECT 107.500000 322.350000 108.500000 323.650000 ;
      RECT 66.500000 322.350000 99.500000 323.650000 ;
      RECT 57.500000 322.350000 58.500000 323.650000 ;
      RECT 29.500000 322.350000 49.500000 323.650000 ;
      RECT 15.500000 322.350000 16.500000 323.650000 ;
      RECT 1157.500000 321.650000 1170.500000 322.350000 ;
      RECT 1107.500000 321.650000 1149.500000 322.350000 ;
      RECT 1057.500000 321.650000 1099.500000 322.350000 ;
      RECT 1007.500000 321.650000 1049.500000 322.350000 ;
      RECT 957.500000 321.650000 999.500000 322.350000 ;
      RECT 907.500000 321.650000 949.500000 322.350000 ;
      RECT 857.500000 321.650000 899.500000 322.350000 ;
      RECT 807.500000 321.650000 849.500000 322.350000 ;
      RECT 757.500000 321.650000 799.500000 322.350000 ;
      RECT 707.500000 321.650000 749.500000 322.350000 ;
      RECT 657.500000 321.650000 699.500000 322.350000 ;
      RECT 607.500000 321.650000 649.500000 322.350000 ;
      RECT 557.500000 321.650000 599.500000 322.350000 ;
      RECT 507.500000 321.650000 549.500000 322.350000 ;
      RECT 457.500000 321.650000 499.500000 322.350000 ;
      RECT 407.500000 321.650000 449.500000 322.350000 ;
      RECT 357.500000 321.650000 399.500000 322.350000 ;
      RECT 307.500000 321.650000 349.500000 322.350000 ;
      RECT 257.500000 321.650000 299.500000 322.350000 ;
      RECT 207.500000 321.650000 249.500000 322.350000 ;
      RECT 157.500000 321.650000 199.500000 322.350000 ;
      RECT 107.500000 321.650000 149.500000 322.350000 ;
      RECT 57.500000 321.650000 99.500000 322.350000 ;
      RECT 15.500000 321.650000 49.500000 322.350000 ;
      RECT 1183.500000 320.350000 1186.000000 323.650000 ;
      RECT 1169.500000 320.350000 1170.500000 321.650000 ;
      RECT 1116.500000 320.350000 1149.500000 321.650000 ;
      RECT 1107.500000 320.350000 1108.500000 321.650000 ;
      RECT 1066.500000 320.350000 1099.500000 321.650000 ;
      RECT 1057.500000 320.350000 1058.500000 321.650000 ;
      RECT 1016.500000 320.350000 1049.500000 321.650000 ;
      RECT 1007.500000 320.350000 1008.500000 321.650000 ;
      RECT 966.500000 320.350000 999.500000 321.650000 ;
      RECT 957.500000 320.350000 958.500000 321.650000 ;
      RECT 916.500000 320.350000 949.500000 321.650000 ;
      RECT 907.500000 320.350000 908.500000 321.650000 ;
      RECT 866.500000 320.350000 899.500000 321.650000 ;
      RECT 857.500000 320.350000 858.500000 321.650000 ;
      RECT 816.500000 320.350000 849.500000 321.650000 ;
      RECT 807.500000 320.350000 808.500000 321.650000 ;
      RECT 766.500000 320.350000 799.500000 321.650000 ;
      RECT 757.500000 320.350000 758.500000 321.650000 ;
      RECT 716.500000 320.350000 749.500000 321.650000 ;
      RECT 707.500000 320.350000 708.500000 321.650000 ;
      RECT 666.500000 320.350000 699.500000 321.650000 ;
      RECT 657.500000 320.350000 658.500000 321.650000 ;
      RECT 616.500000 320.350000 649.500000 321.650000 ;
      RECT 607.500000 320.350000 608.500000 321.650000 ;
      RECT 566.500000 320.350000 599.500000 321.650000 ;
      RECT 557.500000 320.350000 558.500000 321.650000 ;
      RECT 516.500000 320.350000 549.500000 321.650000 ;
      RECT 507.500000 320.350000 508.500000 321.650000 ;
      RECT 466.500000 320.350000 499.500000 321.650000 ;
      RECT 457.500000 320.350000 458.500000 321.650000 ;
      RECT 416.500000 320.350000 449.500000 321.650000 ;
      RECT 407.500000 320.350000 408.500000 321.650000 ;
      RECT 366.500000 320.350000 399.500000 321.650000 ;
      RECT 357.500000 320.350000 358.500000 321.650000 ;
      RECT 316.500000 320.350000 349.500000 321.650000 ;
      RECT 307.500000 320.350000 308.500000 321.650000 ;
      RECT 266.500000 320.350000 299.500000 321.650000 ;
      RECT 257.500000 320.350000 258.500000 321.650000 ;
      RECT 216.500000 320.350000 249.500000 321.650000 ;
      RECT 207.500000 320.350000 208.500000 321.650000 ;
      RECT 166.500000 320.350000 199.500000 321.650000 ;
      RECT 157.500000 320.350000 158.500000 321.650000 ;
      RECT 116.500000 320.350000 149.500000 321.650000 ;
      RECT 107.500000 320.350000 108.500000 321.650000 ;
      RECT 66.500000 320.350000 99.500000 321.650000 ;
      RECT 57.500000 320.350000 58.500000 321.650000 ;
      RECT 29.500000 320.350000 49.500000 321.650000 ;
      RECT 15.500000 320.350000 16.500000 321.650000 ;
      RECT 0.000000 320.350000 2.500000 323.650000 ;
      RECT 1169.500000 319.650000 1186.000000 320.350000 ;
      RECT 1116.500000 319.650000 1156.500000 320.350000 ;
      RECT 1066.500000 319.650000 1108.500000 320.350000 ;
      RECT 1016.500000 319.650000 1058.500000 320.350000 ;
      RECT 966.500000 319.650000 1008.500000 320.350000 ;
      RECT 916.500000 319.650000 958.500000 320.350000 ;
      RECT 866.500000 319.650000 908.500000 320.350000 ;
      RECT 816.500000 319.650000 858.500000 320.350000 ;
      RECT 766.500000 319.650000 808.500000 320.350000 ;
      RECT 716.500000 319.650000 758.500000 320.350000 ;
      RECT 666.500000 319.650000 708.500000 320.350000 ;
      RECT 616.500000 319.650000 658.500000 320.350000 ;
      RECT 566.500000 319.650000 608.500000 320.350000 ;
      RECT 516.500000 319.650000 558.500000 320.350000 ;
      RECT 466.500000 319.650000 508.500000 320.350000 ;
      RECT 366.500000 319.650000 408.500000 320.350000 ;
      RECT 316.500000 319.650000 358.500000 320.350000 ;
      RECT 266.500000 319.650000 308.500000 320.350000 ;
      RECT 216.500000 319.650000 258.500000 320.350000 ;
      RECT 166.500000 319.650000 208.500000 320.350000 ;
      RECT 116.500000 319.650000 158.500000 320.350000 ;
      RECT 66.500000 319.650000 108.500000 320.350000 ;
      RECT 29.500000 319.650000 58.500000 320.350000 ;
      RECT 0.000000 319.650000 16.500000 320.350000 ;
      RECT 416.500000 318.605000 458.500000 320.350000 ;
      RECT 1169.500000 318.350000 1170.500000 319.650000 ;
      RECT 1116.500000 318.350000 1149.500000 319.650000 ;
      RECT 1107.500000 318.350000 1108.500000 319.650000 ;
      RECT 1066.500000 318.350000 1099.500000 319.650000 ;
      RECT 1057.500000 318.350000 1058.500000 319.650000 ;
      RECT 1016.500000 318.350000 1049.500000 319.650000 ;
      RECT 1007.500000 318.350000 1008.500000 319.650000 ;
      RECT 966.500000 318.350000 999.500000 319.650000 ;
      RECT 957.500000 318.350000 958.500000 319.650000 ;
      RECT 916.500000 318.350000 949.500000 319.650000 ;
      RECT 907.500000 318.350000 908.500000 319.650000 ;
      RECT 866.500000 318.350000 899.500000 319.650000 ;
      RECT 857.500000 318.350000 858.500000 319.650000 ;
      RECT 816.500000 318.350000 849.500000 319.650000 ;
      RECT 807.500000 318.350000 808.500000 319.650000 ;
      RECT 766.500000 318.350000 799.500000 319.650000 ;
      RECT 757.500000 318.350000 758.500000 319.650000 ;
      RECT 716.500000 318.350000 749.500000 319.650000 ;
      RECT 707.500000 318.350000 708.500000 319.650000 ;
      RECT 666.500000 318.350000 699.500000 319.650000 ;
      RECT 657.500000 318.350000 658.500000 319.650000 ;
      RECT 616.500000 318.350000 649.500000 319.650000 ;
      RECT 607.500000 318.350000 608.500000 319.650000 ;
      RECT 566.500000 318.350000 599.500000 319.650000 ;
      RECT 557.500000 318.350000 558.500000 319.650000 ;
      RECT 516.500000 318.350000 549.500000 319.650000 ;
      RECT 507.500000 318.350000 508.500000 319.650000 ;
      RECT 466.500000 318.350000 499.500000 319.650000 ;
      RECT 457.500000 318.350000 458.500000 318.605000 ;
      RECT 416.500000 318.350000 449.500000 318.605000 ;
      RECT 407.500000 318.350000 408.500000 319.650000 ;
      RECT 366.500000 318.350000 399.500000 319.650000 ;
      RECT 357.500000 318.350000 358.500000 319.650000 ;
      RECT 316.500000 318.350000 349.500000 319.650000 ;
      RECT 307.500000 318.350000 308.500000 319.650000 ;
      RECT 266.500000 318.350000 299.500000 319.650000 ;
      RECT 257.500000 318.350000 258.500000 319.650000 ;
      RECT 216.500000 318.350000 249.500000 319.650000 ;
      RECT 207.500000 318.350000 208.500000 319.650000 ;
      RECT 166.500000 318.350000 199.500000 319.650000 ;
      RECT 157.500000 318.350000 158.500000 319.650000 ;
      RECT 116.500000 318.350000 149.500000 319.650000 ;
      RECT 107.500000 318.350000 108.500000 319.650000 ;
      RECT 66.500000 318.350000 99.500000 319.650000 ;
      RECT 57.500000 318.350000 58.500000 319.650000 ;
      RECT 29.500000 318.350000 49.500000 319.650000 ;
      RECT 15.500000 318.350000 16.500000 319.650000 ;
      RECT 1157.500000 317.650000 1170.500000 318.350000 ;
      RECT 1107.500000 317.650000 1149.500000 318.350000 ;
      RECT 1057.500000 317.650000 1099.500000 318.350000 ;
      RECT 1007.500000 317.650000 1049.500000 318.350000 ;
      RECT 957.500000 317.650000 999.500000 318.350000 ;
      RECT 907.500000 317.650000 949.500000 318.350000 ;
      RECT 857.500000 317.650000 899.500000 318.350000 ;
      RECT 807.500000 317.650000 849.500000 318.350000 ;
      RECT 757.500000 317.650000 799.500000 318.350000 ;
      RECT 707.500000 317.650000 749.500000 318.350000 ;
      RECT 657.500000 317.650000 699.500000 318.350000 ;
      RECT 607.500000 317.650000 649.500000 318.350000 ;
      RECT 557.500000 317.650000 599.500000 318.350000 ;
      RECT 507.500000 317.650000 549.500000 318.350000 ;
      RECT 407.500000 317.650000 449.500000 318.350000 ;
      RECT 357.500000 317.650000 399.500000 318.350000 ;
      RECT 307.500000 317.650000 349.500000 318.350000 ;
      RECT 257.500000 317.650000 299.500000 318.350000 ;
      RECT 207.500000 317.650000 249.500000 318.350000 ;
      RECT 157.500000 317.650000 199.500000 318.350000 ;
      RECT 107.500000 317.650000 149.500000 318.350000 ;
      RECT 57.500000 317.650000 99.500000 318.350000 ;
      RECT 15.500000 317.650000 49.500000 318.350000 ;
      RECT 1183.500000 316.350000 1186.000000 319.650000 ;
      RECT 1169.500000 316.350000 1170.500000 317.650000 ;
      RECT 1116.500000 316.350000 1149.500000 317.650000 ;
      RECT 1107.500000 316.350000 1108.500000 317.650000 ;
      RECT 1066.500000 316.350000 1099.500000 317.650000 ;
      RECT 1057.500000 316.350000 1058.500000 317.650000 ;
      RECT 1016.500000 316.350000 1049.500000 317.650000 ;
      RECT 1007.500000 316.350000 1008.500000 317.650000 ;
      RECT 966.500000 316.350000 999.500000 317.650000 ;
      RECT 957.500000 316.350000 958.500000 317.650000 ;
      RECT 916.500000 316.350000 949.500000 317.650000 ;
      RECT 907.500000 316.350000 908.500000 317.650000 ;
      RECT 866.500000 316.350000 899.500000 317.650000 ;
      RECT 857.500000 316.350000 858.500000 317.650000 ;
      RECT 816.500000 316.350000 849.500000 317.650000 ;
      RECT 807.500000 316.350000 808.500000 317.650000 ;
      RECT 766.500000 316.350000 799.500000 317.650000 ;
      RECT 757.500000 316.350000 758.500000 317.650000 ;
      RECT 716.500000 316.350000 749.500000 317.650000 ;
      RECT 707.500000 316.350000 708.500000 317.650000 ;
      RECT 666.500000 316.350000 699.500000 317.650000 ;
      RECT 657.500000 316.350000 658.500000 317.650000 ;
      RECT 616.500000 316.350000 649.500000 317.650000 ;
      RECT 607.500000 316.350000 608.500000 317.650000 ;
      RECT 566.500000 316.350000 599.500000 317.650000 ;
      RECT 557.500000 316.350000 558.500000 317.650000 ;
      RECT 516.500000 316.350000 549.500000 317.650000 ;
      RECT 507.500000 316.350000 508.500000 317.650000 ;
      RECT 457.500000 316.350000 499.500000 318.350000 ;
      RECT 407.500000 316.350000 408.500000 317.650000 ;
      RECT 366.500000 316.350000 399.500000 317.650000 ;
      RECT 357.500000 316.350000 358.500000 317.650000 ;
      RECT 316.500000 316.350000 349.500000 317.650000 ;
      RECT 307.500000 316.350000 308.500000 317.650000 ;
      RECT 266.500000 316.350000 299.500000 317.650000 ;
      RECT 257.500000 316.350000 258.500000 317.650000 ;
      RECT 216.500000 316.350000 249.500000 317.650000 ;
      RECT 207.500000 316.350000 208.500000 317.650000 ;
      RECT 166.500000 316.350000 199.500000 317.650000 ;
      RECT 157.500000 316.350000 158.500000 317.650000 ;
      RECT 116.500000 316.350000 149.500000 317.650000 ;
      RECT 107.500000 316.350000 108.500000 317.650000 ;
      RECT 66.500000 316.350000 99.500000 317.650000 ;
      RECT 57.500000 316.350000 58.500000 317.650000 ;
      RECT 29.500000 316.350000 49.500000 317.650000 ;
      RECT 15.500000 316.350000 16.500000 317.650000 ;
      RECT 0.000000 316.350000 2.500000 319.650000 ;
      RECT 1169.500000 315.650000 1186.000000 316.350000 ;
      RECT 1116.500000 315.650000 1156.500000 316.350000 ;
      RECT 1066.500000 315.650000 1108.500000 316.350000 ;
      RECT 1016.500000 315.650000 1058.500000 316.350000 ;
      RECT 966.500000 315.650000 1008.500000 316.350000 ;
      RECT 916.500000 315.650000 958.500000 316.350000 ;
      RECT 866.500000 315.650000 908.500000 316.350000 ;
      RECT 816.500000 315.650000 858.500000 316.350000 ;
      RECT 766.500000 315.650000 808.500000 316.350000 ;
      RECT 716.500000 315.650000 758.500000 316.350000 ;
      RECT 666.500000 315.650000 708.500000 316.350000 ;
      RECT 616.500000 315.650000 658.500000 316.350000 ;
      RECT 566.500000 315.650000 608.500000 316.350000 ;
      RECT 516.500000 315.650000 558.500000 316.350000 ;
      RECT 457.500000 315.650000 508.500000 316.350000 ;
      RECT 366.500000 315.650000 408.500000 316.350000 ;
      RECT 316.500000 315.650000 358.500000 316.350000 ;
      RECT 266.500000 315.650000 308.500000 316.350000 ;
      RECT 216.500000 315.650000 258.500000 316.350000 ;
      RECT 166.500000 315.650000 208.500000 316.350000 ;
      RECT 116.500000 315.650000 158.500000 316.350000 ;
      RECT 66.500000 315.650000 108.500000 316.350000 ;
      RECT 29.500000 315.650000 58.500000 316.350000 ;
      RECT 0.000000 315.650000 16.500000 316.350000 ;
      RECT 457.500000 314.605000 499.500000 315.650000 ;
      RECT 416.500000 314.605000 449.500000 317.650000 ;
      RECT 1169.500000 314.350000 1170.500000 315.650000 ;
      RECT 1116.500000 314.350000 1149.500000 315.650000 ;
      RECT 1107.500000 314.350000 1108.500000 315.650000 ;
      RECT 1066.500000 314.350000 1099.500000 315.650000 ;
      RECT 1057.500000 314.350000 1058.500000 315.650000 ;
      RECT 1016.500000 314.350000 1049.500000 315.650000 ;
      RECT 1007.500000 314.350000 1008.500000 315.650000 ;
      RECT 966.500000 314.350000 999.500000 315.650000 ;
      RECT 957.500000 314.350000 958.500000 315.650000 ;
      RECT 916.500000 314.350000 949.500000 315.650000 ;
      RECT 907.500000 314.350000 908.500000 315.650000 ;
      RECT 866.500000 314.350000 899.500000 315.650000 ;
      RECT 857.500000 314.350000 858.500000 315.650000 ;
      RECT 816.500000 314.350000 849.500000 315.650000 ;
      RECT 807.500000 314.350000 808.500000 315.650000 ;
      RECT 766.500000 314.350000 799.500000 315.650000 ;
      RECT 757.500000 314.350000 758.500000 315.650000 ;
      RECT 716.500000 314.350000 749.500000 315.650000 ;
      RECT 707.500000 314.350000 708.500000 315.650000 ;
      RECT 666.500000 314.350000 699.500000 315.650000 ;
      RECT 657.500000 314.350000 658.500000 315.650000 ;
      RECT 616.500000 314.350000 649.500000 315.650000 ;
      RECT 607.500000 314.350000 608.500000 315.650000 ;
      RECT 566.500000 314.350000 599.500000 315.650000 ;
      RECT 557.500000 314.350000 558.500000 315.650000 ;
      RECT 516.500000 314.350000 549.500000 315.650000 ;
      RECT 507.500000 314.350000 508.500000 315.650000 ;
      RECT 416.500000 314.350000 499.500000 314.605000 ;
      RECT 407.500000 314.350000 408.500000 315.650000 ;
      RECT 366.500000 314.350000 399.500000 315.650000 ;
      RECT 357.500000 314.350000 358.500000 315.650000 ;
      RECT 316.500000 314.350000 349.500000 315.650000 ;
      RECT 307.500000 314.350000 308.500000 315.650000 ;
      RECT 266.500000 314.350000 299.500000 315.650000 ;
      RECT 257.500000 314.350000 258.500000 315.650000 ;
      RECT 216.500000 314.350000 249.500000 315.650000 ;
      RECT 207.500000 314.350000 208.500000 315.650000 ;
      RECT 166.500000 314.350000 199.500000 315.650000 ;
      RECT 157.500000 314.350000 158.500000 315.650000 ;
      RECT 116.500000 314.350000 149.500000 315.650000 ;
      RECT 107.500000 314.350000 108.500000 315.650000 ;
      RECT 66.500000 314.350000 99.500000 315.650000 ;
      RECT 57.500000 314.350000 58.500000 315.650000 ;
      RECT 29.500000 314.350000 49.500000 315.650000 ;
      RECT 15.500000 314.350000 16.500000 315.650000 ;
      RECT 1157.500000 313.650000 1170.500000 314.350000 ;
      RECT 1107.500000 313.650000 1149.500000 314.350000 ;
      RECT 1057.500000 313.650000 1099.500000 314.350000 ;
      RECT 1007.500000 313.650000 1049.500000 314.350000 ;
      RECT 957.500000 313.650000 999.500000 314.350000 ;
      RECT 907.500000 313.650000 949.500000 314.350000 ;
      RECT 857.500000 313.650000 899.500000 314.350000 ;
      RECT 807.500000 313.650000 849.500000 314.350000 ;
      RECT 757.500000 313.650000 799.500000 314.350000 ;
      RECT 707.500000 313.650000 749.500000 314.350000 ;
      RECT 657.500000 313.650000 699.500000 314.350000 ;
      RECT 607.500000 313.650000 649.500000 314.350000 ;
      RECT 557.500000 313.650000 599.500000 314.350000 ;
      RECT 507.500000 313.650000 549.500000 314.350000 ;
      RECT 407.500000 313.650000 499.500000 314.350000 ;
      RECT 357.500000 313.650000 399.500000 314.350000 ;
      RECT 307.500000 313.650000 349.500000 314.350000 ;
      RECT 257.500000 313.650000 299.500000 314.350000 ;
      RECT 207.500000 313.650000 249.500000 314.350000 ;
      RECT 157.500000 313.650000 199.500000 314.350000 ;
      RECT 107.500000 313.650000 149.500000 314.350000 ;
      RECT 57.500000 313.650000 99.500000 314.350000 ;
      RECT 15.500000 313.650000 49.500000 314.350000 ;
      RECT 1183.500000 312.350000 1186.000000 315.650000 ;
      RECT 1169.500000 312.350000 1170.500000 313.650000 ;
      RECT 1116.500000 312.350000 1149.500000 313.650000 ;
      RECT 1107.500000 312.350000 1108.500000 313.650000 ;
      RECT 1066.500000 312.350000 1099.500000 313.650000 ;
      RECT 1057.500000 312.350000 1058.500000 313.650000 ;
      RECT 1016.500000 312.350000 1049.500000 313.650000 ;
      RECT 1007.500000 312.350000 1008.500000 313.650000 ;
      RECT 966.500000 312.350000 999.500000 313.650000 ;
      RECT 957.500000 312.350000 958.500000 313.650000 ;
      RECT 916.500000 312.350000 949.500000 313.650000 ;
      RECT 907.500000 312.350000 908.500000 313.650000 ;
      RECT 866.500000 312.350000 899.500000 313.650000 ;
      RECT 857.500000 312.350000 858.500000 313.650000 ;
      RECT 816.500000 312.350000 849.500000 313.650000 ;
      RECT 807.500000 312.350000 808.500000 313.650000 ;
      RECT 766.500000 312.350000 799.500000 313.650000 ;
      RECT 757.500000 312.350000 758.500000 313.650000 ;
      RECT 716.500000 312.350000 749.500000 313.650000 ;
      RECT 707.500000 312.350000 708.500000 313.650000 ;
      RECT 666.500000 312.350000 699.500000 313.650000 ;
      RECT 657.500000 312.350000 658.500000 313.650000 ;
      RECT 616.500000 312.350000 649.500000 313.650000 ;
      RECT 607.500000 312.350000 608.500000 313.650000 ;
      RECT 566.500000 312.350000 599.500000 313.650000 ;
      RECT 557.500000 312.350000 558.500000 313.650000 ;
      RECT 516.500000 312.350000 549.500000 313.650000 ;
      RECT 507.500000 312.350000 508.500000 313.650000 ;
      RECT 416.500000 312.350000 499.500000 313.650000 ;
      RECT 407.500000 312.350000 408.500000 313.650000 ;
      RECT 366.500000 312.350000 399.500000 313.650000 ;
      RECT 357.500000 312.350000 358.500000 313.650000 ;
      RECT 316.500000 312.350000 349.500000 313.650000 ;
      RECT 307.500000 312.350000 308.500000 313.650000 ;
      RECT 266.500000 312.350000 299.500000 313.650000 ;
      RECT 257.500000 312.350000 258.500000 313.650000 ;
      RECT 216.500000 312.350000 249.500000 313.650000 ;
      RECT 207.500000 312.350000 208.500000 313.650000 ;
      RECT 166.500000 312.350000 199.500000 313.650000 ;
      RECT 157.500000 312.350000 158.500000 313.650000 ;
      RECT 116.500000 312.350000 149.500000 313.650000 ;
      RECT 107.500000 312.350000 108.500000 313.650000 ;
      RECT 66.500000 312.350000 99.500000 313.650000 ;
      RECT 57.500000 312.350000 58.500000 313.650000 ;
      RECT 29.500000 312.350000 49.500000 313.650000 ;
      RECT 15.500000 312.350000 16.500000 313.650000 ;
      RECT 0.000000 312.350000 2.500000 315.650000 ;
      RECT 1169.500000 311.650000 1186.000000 312.350000 ;
      RECT 1116.500000 311.650000 1156.500000 312.350000 ;
      RECT 1066.500000 311.650000 1108.500000 312.350000 ;
      RECT 1016.500000 311.650000 1058.500000 312.350000 ;
      RECT 966.500000 311.650000 1008.500000 312.350000 ;
      RECT 916.500000 311.650000 958.500000 312.350000 ;
      RECT 866.500000 311.650000 908.500000 312.350000 ;
      RECT 816.500000 311.650000 858.500000 312.350000 ;
      RECT 766.500000 311.650000 808.500000 312.350000 ;
      RECT 716.500000 311.650000 758.500000 312.350000 ;
      RECT 666.500000 311.650000 708.500000 312.350000 ;
      RECT 616.500000 311.650000 658.500000 312.350000 ;
      RECT 566.500000 311.650000 608.500000 312.350000 ;
      RECT 516.500000 311.650000 558.500000 312.350000 ;
      RECT 416.500000 311.650000 508.500000 312.350000 ;
      RECT 366.500000 311.650000 408.500000 312.350000 ;
      RECT 316.500000 311.650000 358.500000 312.350000 ;
      RECT 266.500000 311.650000 308.500000 312.350000 ;
      RECT 216.500000 311.650000 258.500000 312.350000 ;
      RECT 166.500000 311.650000 208.500000 312.350000 ;
      RECT 116.500000 311.650000 158.500000 312.350000 ;
      RECT 66.500000 311.650000 108.500000 312.350000 ;
      RECT 29.500000 311.650000 58.500000 312.350000 ;
      RECT 0.000000 311.650000 16.500000 312.350000 ;
      RECT 1169.500000 310.350000 1170.500000 311.650000 ;
      RECT 1116.500000 310.350000 1149.500000 311.650000 ;
      RECT 1107.500000 310.350000 1108.500000 311.650000 ;
      RECT 1066.500000 310.350000 1099.500000 311.650000 ;
      RECT 1057.500000 310.350000 1058.500000 311.650000 ;
      RECT 1016.500000 310.350000 1049.500000 311.650000 ;
      RECT 1007.500000 310.350000 1008.500000 311.650000 ;
      RECT 966.500000 310.350000 999.500000 311.650000 ;
      RECT 957.500000 310.350000 958.500000 311.650000 ;
      RECT 916.500000 310.350000 949.500000 311.650000 ;
      RECT 907.500000 310.350000 908.500000 311.650000 ;
      RECT 866.500000 310.350000 899.500000 311.650000 ;
      RECT 857.500000 310.350000 858.500000 311.650000 ;
      RECT 816.500000 310.350000 849.500000 311.650000 ;
      RECT 807.500000 310.350000 808.500000 311.650000 ;
      RECT 766.500000 310.350000 799.500000 311.650000 ;
      RECT 757.500000 310.350000 758.500000 311.650000 ;
      RECT 716.500000 310.350000 749.500000 311.650000 ;
      RECT 707.500000 310.350000 708.500000 311.650000 ;
      RECT 666.500000 310.350000 699.500000 311.650000 ;
      RECT 657.500000 310.350000 658.500000 311.650000 ;
      RECT 616.500000 310.350000 649.500000 311.650000 ;
      RECT 607.500000 310.350000 608.500000 311.650000 ;
      RECT 566.500000 310.350000 599.500000 311.650000 ;
      RECT 557.500000 310.350000 558.500000 311.650000 ;
      RECT 516.500000 310.350000 549.500000 311.650000 ;
      RECT 507.500000 310.350000 508.500000 311.650000 ;
      RECT 416.500000 310.350000 499.500000 311.650000 ;
      RECT 407.500000 310.350000 408.500000 311.650000 ;
      RECT 366.500000 310.350000 399.500000 311.650000 ;
      RECT 357.500000 310.350000 358.500000 311.650000 ;
      RECT 316.500000 310.350000 349.500000 311.650000 ;
      RECT 307.500000 310.350000 308.500000 311.650000 ;
      RECT 266.500000 310.350000 299.500000 311.650000 ;
      RECT 257.500000 310.350000 258.500000 311.650000 ;
      RECT 216.500000 310.350000 249.500000 311.650000 ;
      RECT 207.500000 310.350000 208.500000 311.650000 ;
      RECT 166.500000 310.350000 199.500000 311.650000 ;
      RECT 157.500000 310.350000 158.500000 311.650000 ;
      RECT 116.500000 310.350000 149.500000 311.650000 ;
      RECT 107.500000 310.350000 108.500000 311.650000 ;
      RECT 66.500000 310.350000 99.500000 311.650000 ;
      RECT 57.500000 310.350000 58.500000 311.650000 ;
      RECT 29.500000 310.350000 49.500000 311.650000 ;
      RECT 15.500000 310.350000 16.500000 311.650000 ;
      RECT 1157.500000 309.650000 1170.500000 310.350000 ;
      RECT 1107.500000 309.650000 1149.500000 310.350000 ;
      RECT 1057.500000 309.650000 1099.500000 310.350000 ;
      RECT 1007.500000 309.650000 1049.500000 310.350000 ;
      RECT 957.500000 309.650000 999.500000 310.350000 ;
      RECT 907.500000 309.650000 949.500000 310.350000 ;
      RECT 857.500000 309.650000 899.500000 310.350000 ;
      RECT 807.500000 309.650000 849.500000 310.350000 ;
      RECT 757.500000 309.650000 799.500000 310.350000 ;
      RECT 707.500000 309.650000 749.500000 310.350000 ;
      RECT 657.500000 309.650000 699.500000 310.350000 ;
      RECT 607.500000 309.650000 649.500000 310.350000 ;
      RECT 557.500000 309.650000 599.500000 310.350000 ;
      RECT 507.500000 309.650000 549.500000 310.350000 ;
      RECT 407.500000 309.650000 499.500000 310.350000 ;
      RECT 357.500000 309.650000 399.500000 310.350000 ;
      RECT 307.500000 309.650000 349.500000 310.350000 ;
      RECT 257.500000 309.650000 299.500000 310.350000 ;
      RECT 207.500000 309.650000 249.500000 310.350000 ;
      RECT 157.500000 309.650000 199.500000 310.350000 ;
      RECT 107.500000 309.650000 149.500000 310.350000 ;
      RECT 57.500000 309.650000 99.500000 310.350000 ;
      RECT 15.500000 309.650000 49.500000 310.350000 ;
      RECT 1183.500000 308.350000 1186.000000 311.650000 ;
      RECT 1169.500000 308.350000 1170.500000 309.650000 ;
      RECT 1116.500000 308.350000 1149.500000 309.650000 ;
      RECT 1107.500000 308.350000 1108.500000 309.650000 ;
      RECT 1066.500000 308.350000 1099.500000 309.650000 ;
      RECT 1057.500000 308.350000 1058.500000 309.650000 ;
      RECT 1016.500000 308.350000 1049.500000 309.650000 ;
      RECT 1007.500000 308.350000 1008.500000 309.650000 ;
      RECT 966.500000 308.350000 999.500000 309.650000 ;
      RECT 957.500000 308.350000 958.500000 309.650000 ;
      RECT 916.500000 308.350000 949.500000 309.650000 ;
      RECT 907.500000 308.350000 908.500000 309.650000 ;
      RECT 866.500000 308.350000 899.500000 309.650000 ;
      RECT 857.500000 308.350000 858.500000 309.650000 ;
      RECT 816.500000 308.350000 849.500000 309.650000 ;
      RECT 807.500000 308.350000 808.500000 309.650000 ;
      RECT 766.500000 308.350000 799.500000 309.650000 ;
      RECT 757.500000 308.350000 758.500000 309.650000 ;
      RECT 716.500000 308.350000 749.500000 309.650000 ;
      RECT 707.500000 308.350000 708.500000 309.650000 ;
      RECT 666.500000 308.350000 699.500000 309.650000 ;
      RECT 657.500000 308.350000 658.500000 309.650000 ;
      RECT 616.500000 308.350000 649.500000 309.650000 ;
      RECT 607.500000 308.350000 608.500000 309.650000 ;
      RECT 566.500000 308.350000 599.500000 309.650000 ;
      RECT 557.500000 308.350000 558.500000 309.650000 ;
      RECT 516.500000 308.350000 549.500000 309.650000 ;
      RECT 507.500000 308.350000 508.500000 309.650000 ;
      RECT 416.500000 308.350000 499.500000 309.650000 ;
      RECT 407.500000 308.350000 408.500000 309.650000 ;
      RECT 366.500000 308.350000 399.500000 309.650000 ;
      RECT 357.500000 308.350000 358.500000 309.650000 ;
      RECT 316.500000 308.350000 349.500000 309.650000 ;
      RECT 307.500000 308.350000 308.500000 309.650000 ;
      RECT 266.500000 308.350000 299.500000 309.650000 ;
      RECT 257.500000 308.350000 258.500000 309.650000 ;
      RECT 216.500000 308.350000 249.500000 309.650000 ;
      RECT 207.500000 308.350000 208.500000 309.650000 ;
      RECT 166.500000 308.350000 199.500000 309.650000 ;
      RECT 157.500000 308.350000 158.500000 309.650000 ;
      RECT 116.500000 308.350000 149.500000 309.650000 ;
      RECT 107.500000 308.350000 108.500000 309.650000 ;
      RECT 66.500000 308.350000 99.500000 309.650000 ;
      RECT 57.500000 308.350000 58.500000 309.650000 ;
      RECT 29.500000 308.350000 49.500000 309.650000 ;
      RECT 15.500000 308.350000 16.500000 309.650000 ;
      RECT 0.000000 308.350000 2.500000 311.650000 ;
      RECT 1169.500000 307.650000 1186.000000 308.350000 ;
      RECT 1116.500000 307.650000 1156.500000 308.350000 ;
      RECT 1066.500000 307.650000 1108.500000 308.350000 ;
      RECT 1016.500000 307.650000 1058.500000 308.350000 ;
      RECT 966.500000 307.650000 1008.500000 308.350000 ;
      RECT 916.500000 307.650000 958.500000 308.350000 ;
      RECT 866.500000 307.650000 908.500000 308.350000 ;
      RECT 816.500000 307.650000 858.500000 308.350000 ;
      RECT 766.500000 307.650000 808.500000 308.350000 ;
      RECT 716.500000 307.650000 758.500000 308.350000 ;
      RECT 666.500000 307.650000 708.500000 308.350000 ;
      RECT 616.500000 307.650000 658.500000 308.350000 ;
      RECT 566.500000 307.650000 608.500000 308.350000 ;
      RECT 516.500000 307.650000 558.500000 308.350000 ;
      RECT 416.500000 307.650000 508.500000 308.350000 ;
      RECT 366.500000 307.650000 408.500000 308.350000 ;
      RECT 316.500000 307.650000 358.500000 308.350000 ;
      RECT 266.500000 307.650000 308.500000 308.350000 ;
      RECT 216.500000 307.650000 258.500000 308.350000 ;
      RECT 166.500000 307.650000 208.500000 308.350000 ;
      RECT 116.500000 307.650000 158.500000 308.350000 ;
      RECT 66.500000 307.650000 108.500000 308.350000 ;
      RECT 29.500000 307.650000 58.500000 308.350000 ;
      RECT 0.000000 307.650000 16.500000 308.350000 ;
      RECT 1169.500000 306.350000 1170.500000 307.650000 ;
      RECT 1116.500000 306.350000 1149.500000 307.650000 ;
      RECT 1107.500000 306.350000 1108.500000 307.650000 ;
      RECT 1066.500000 306.350000 1099.500000 307.650000 ;
      RECT 1057.500000 306.350000 1058.500000 307.650000 ;
      RECT 1016.500000 306.350000 1049.500000 307.650000 ;
      RECT 1007.500000 306.350000 1008.500000 307.650000 ;
      RECT 966.500000 306.350000 999.500000 307.650000 ;
      RECT 957.500000 306.350000 958.500000 307.650000 ;
      RECT 916.500000 306.350000 949.500000 307.650000 ;
      RECT 907.500000 306.350000 908.500000 307.650000 ;
      RECT 866.500000 306.350000 899.500000 307.650000 ;
      RECT 857.500000 306.350000 858.500000 307.650000 ;
      RECT 816.500000 306.350000 849.500000 307.650000 ;
      RECT 807.500000 306.350000 808.500000 307.650000 ;
      RECT 766.500000 306.350000 799.500000 307.650000 ;
      RECT 757.500000 306.350000 758.500000 307.650000 ;
      RECT 716.500000 306.350000 749.500000 307.650000 ;
      RECT 707.500000 306.350000 708.500000 307.650000 ;
      RECT 666.500000 306.350000 699.500000 307.650000 ;
      RECT 657.500000 306.350000 658.500000 307.650000 ;
      RECT 616.500000 306.350000 649.500000 307.650000 ;
      RECT 607.500000 306.350000 608.500000 307.650000 ;
      RECT 566.500000 306.350000 599.500000 307.650000 ;
      RECT 557.500000 306.350000 558.500000 307.650000 ;
      RECT 516.500000 306.350000 549.500000 307.650000 ;
      RECT 507.500000 306.350000 508.500000 307.650000 ;
      RECT 416.500000 306.350000 499.500000 307.650000 ;
      RECT 407.500000 306.350000 408.500000 307.650000 ;
      RECT 366.500000 306.350000 399.500000 307.650000 ;
      RECT 357.500000 306.350000 358.500000 307.650000 ;
      RECT 316.500000 306.350000 349.500000 307.650000 ;
      RECT 307.500000 306.350000 308.500000 307.650000 ;
      RECT 266.500000 306.350000 299.500000 307.650000 ;
      RECT 257.500000 306.350000 258.500000 307.650000 ;
      RECT 216.500000 306.350000 249.500000 307.650000 ;
      RECT 207.500000 306.350000 208.500000 307.650000 ;
      RECT 166.500000 306.350000 199.500000 307.650000 ;
      RECT 157.500000 306.350000 158.500000 307.650000 ;
      RECT 116.500000 306.350000 149.500000 307.650000 ;
      RECT 107.500000 306.350000 108.500000 307.650000 ;
      RECT 66.500000 306.350000 99.500000 307.650000 ;
      RECT 57.500000 306.350000 58.500000 307.650000 ;
      RECT 29.500000 306.350000 49.500000 307.650000 ;
      RECT 15.500000 306.350000 16.500000 307.650000 ;
      RECT 1157.500000 305.650000 1170.500000 306.350000 ;
      RECT 1107.500000 305.650000 1149.500000 306.350000 ;
      RECT 1057.500000 305.650000 1099.500000 306.350000 ;
      RECT 1007.500000 305.650000 1049.500000 306.350000 ;
      RECT 957.500000 305.650000 999.500000 306.350000 ;
      RECT 907.500000 305.650000 949.500000 306.350000 ;
      RECT 857.500000 305.650000 899.500000 306.350000 ;
      RECT 807.500000 305.650000 849.500000 306.350000 ;
      RECT 757.500000 305.650000 799.500000 306.350000 ;
      RECT 707.500000 305.650000 749.500000 306.350000 ;
      RECT 657.500000 305.650000 699.500000 306.350000 ;
      RECT 607.500000 305.650000 649.500000 306.350000 ;
      RECT 557.500000 305.650000 599.500000 306.350000 ;
      RECT 507.500000 305.650000 549.500000 306.350000 ;
      RECT 407.500000 305.650000 499.500000 306.350000 ;
      RECT 357.500000 305.650000 399.500000 306.350000 ;
      RECT 307.500000 305.650000 349.500000 306.350000 ;
      RECT 257.500000 305.650000 299.500000 306.350000 ;
      RECT 207.500000 305.650000 249.500000 306.350000 ;
      RECT 157.500000 305.650000 199.500000 306.350000 ;
      RECT 107.500000 305.650000 149.500000 306.350000 ;
      RECT 57.500000 305.650000 99.500000 306.350000 ;
      RECT 15.500000 305.650000 49.500000 306.350000 ;
      RECT 1183.500000 304.350000 1186.000000 307.650000 ;
      RECT 1169.500000 304.350000 1170.500000 305.650000 ;
      RECT 1116.500000 304.350000 1149.500000 305.650000 ;
      RECT 1107.500000 304.350000 1108.500000 305.650000 ;
      RECT 1066.500000 304.350000 1099.500000 305.650000 ;
      RECT 1057.500000 304.350000 1058.500000 305.650000 ;
      RECT 1016.500000 304.350000 1049.500000 305.650000 ;
      RECT 1007.500000 304.350000 1008.500000 305.650000 ;
      RECT 966.500000 304.350000 999.500000 305.650000 ;
      RECT 957.500000 304.350000 958.500000 305.650000 ;
      RECT 916.500000 304.350000 949.500000 305.650000 ;
      RECT 907.500000 304.350000 908.500000 305.650000 ;
      RECT 866.500000 304.350000 899.500000 305.650000 ;
      RECT 857.500000 304.350000 858.500000 305.650000 ;
      RECT 816.500000 304.350000 849.500000 305.650000 ;
      RECT 807.500000 304.350000 808.500000 305.650000 ;
      RECT 766.500000 304.350000 799.500000 305.650000 ;
      RECT 757.500000 304.350000 758.500000 305.650000 ;
      RECT 716.500000 304.350000 749.500000 305.650000 ;
      RECT 707.500000 304.350000 708.500000 305.650000 ;
      RECT 666.500000 304.350000 699.500000 305.650000 ;
      RECT 657.500000 304.350000 658.500000 305.650000 ;
      RECT 616.500000 304.350000 649.500000 305.650000 ;
      RECT 607.500000 304.350000 608.500000 305.650000 ;
      RECT 566.500000 304.350000 599.500000 305.650000 ;
      RECT 557.500000 304.350000 558.500000 305.650000 ;
      RECT 516.500000 304.350000 549.500000 305.650000 ;
      RECT 507.500000 304.350000 508.500000 305.650000 ;
      RECT 416.500000 304.350000 499.500000 305.650000 ;
      RECT 407.500000 304.350000 408.500000 305.650000 ;
      RECT 366.500000 304.350000 399.500000 305.650000 ;
      RECT 357.500000 304.350000 358.500000 305.650000 ;
      RECT 316.500000 304.350000 349.500000 305.650000 ;
      RECT 307.500000 304.350000 308.500000 305.650000 ;
      RECT 266.500000 304.350000 299.500000 305.650000 ;
      RECT 257.500000 304.350000 258.500000 305.650000 ;
      RECT 216.500000 304.350000 249.500000 305.650000 ;
      RECT 207.500000 304.350000 208.500000 305.650000 ;
      RECT 166.500000 304.350000 199.500000 305.650000 ;
      RECT 157.500000 304.350000 158.500000 305.650000 ;
      RECT 116.500000 304.350000 149.500000 305.650000 ;
      RECT 107.500000 304.350000 108.500000 305.650000 ;
      RECT 66.500000 304.350000 99.500000 305.650000 ;
      RECT 57.500000 304.350000 58.500000 305.650000 ;
      RECT 29.500000 304.350000 49.500000 305.650000 ;
      RECT 15.500000 304.350000 16.500000 305.650000 ;
      RECT 0.000000 304.350000 2.500000 307.650000 ;
      RECT 416.500000 303.730000 508.500000 304.350000 ;
      RECT 1169.500000 303.650000 1186.000000 304.350000 ;
      RECT 1116.500000 303.650000 1156.500000 304.350000 ;
      RECT 1066.500000 303.650000 1108.500000 304.350000 ;
      RECT 1016.500000 303.650000 1058.500000 304.350000 ;
      RECT 966.500000 303.650000 1008.500000 304.350000 ;
      RECT 916.500000 303.650000 958.500000 304.350000 ;
      RECT 866.500000 303.650000 908.500000 304.350000 ;
      RECT 816.500000 303.650000 858.500000 304.350000 ;
      RECT 766.500000 303.650000 808.500000 304.350000 ;
      RECT 716.500000 303.650000 758.500000 304.350000 ;
      RECT 666.500000 303.650000 708.500000 304.350000 ;
      RECT 616.500000 303.650000 658.500000 304.350000 ;
      RECT 566.500000 303.650000 608.500000 304.350000 ;
      RECT 516.500000 303.650000 558.500000 304.350000 ;
      RECT 466.500000 303.650000 508.500000 303.730000 ;
      RECT 366.500000 303.650000 408.500000 304.350000 ;
      RECT 316.500000 303.650000 358.500000 304.350000 ;
      RECT 266.500000 303.650000 308.500000 304.350000 ;
      RECT 216.500000 303.650000 258.500000 304.350000 ;
      RECT 166.500000 303.650000 208.500000 304.350000 ;
      RECT 116.500000 303.650000 158.500000 304.350000 ;
      RECT 66.500000 303.650000 108.500000 304.350000 ;
      RECT 29.500000 303.650000 58.500000 304.350000 ;
      RECT 0.000000 303.650000 16.500000 304.350000 ;
      RECT 1169.500000 302.350000 1170.500000 303.650000 ;
      RECT 1116.500000 302.350000 1149.500000 303.650000 ;
      RECT 1107.500000 302.350000 1108.500000 303.650000 ;
      RECT 1066.500000 302.350000 1099.500000 303.650000 ;
      RECT 1057.500000 302.350000 1058.500000 303.650000 ;
      RECT 1016.500000 302.350000 1049.500000 303.650000 ;
      RECT 1007.500000 302.350000 1008.500000 303.650000 ;
      RECT 966.500000 302.350000 999.500000 303.650000 ;
      RECT 957.500000 302.350000 958.500000 303.650000 ;
      RECT 916.500000 302.350000 949.500000 303.650000 ;
      RECT 907.500000 302.350000 908.500000 303.650000 ;
      RECT 866.500000 302.350000 899.500000 303.650000 ;
      RECT 857.500000 302.350000 858.500000 303.650000 ;
      RECT 816.500000 302.350000 849.500000 303.650000 ;
      RECT 807.500000 302.350000 808.500000 303.650000 ;
      RECT 766.500000 302.350000 799.500000 303.650000 ;
      RECT 757.500000 302.350000 758.500000 303.650000 ;
      RECT 716.500000 302.350000 749.500000 303.650000 ;
      RECT 707.500000 302.350000 708.500000 303.650000 ;
      RECT 666.500000 302.350000 699.500000 303.650000 ;
      RECT 657.500000 302.350000 658.500000 303.650000 ;
      RECT 616.500000 302.350000 649.500000 303.650000 ;
      RECT 607.500000 302.350000 608.500000 303.650000 ;
      RECT 566.500000 302.350000 599.500000 303.650000 ;
      RECT 557.500000 302.350000 558.500000 303.650000 ;
      RECT 516.500000 302.350000 549.500000 303.650000 ;
      RECT 507.500000 302.350000 508.500000 303.650000 ;
      RECT 416.500000 302.350000 458.500000 303.730000 ;
      RECT 407.500000 302.350000 408.500000 303.650000 ;
      RECT 366.500000 302.350000 399.500000 303.650000 ;
      RECT 357.500000 302.350000 358.500000 303.650000 ;
      RECT 316.500000 302.350000 349.500000 303.650000 ;
      RECT 307.500000 302.350000 308.500000 303.650000 ;
      RECT 266.500000 302.350000 299.500000 303.650000 ;
      RECT 257.500000 302.350000 258.500000 303.650000 ;
      RECT 216.500000 302.350000 249.500000 303.650000 ;
      RECT 207.500000 302.350000 208.500000 303.650000 ;
      RECT 166.500000 302.350000 199.500000 303.650000 ;
      RECT 157.500000 302.350000 158.500000 303.650000 ;
      RECT 116.500000 302.350000 149.500000 303.650000 ;
      RECT 107.500000 302.350000 108.500000 303.650000 ;
      RECT 66.500000 302.350000 99.500000 303.650000 ;
      RECT 57.500000 302.350000 58.500000 303.650000 ;
      RECT 29.500000 302.350000 49.500000 303.650000 ;
      RECT 15.500000 302.350000 16.500000 303.650000 ;
      RECT 1157.500000 301.650000 1170.500000 302.350000 ;
      RECT 1107.500000 301.650000 1149.500000 302.350000 ;
      RECT 1057.500000 301.650000 1099.500000 302.350000 ;
      RECT 1007.500000 301.650000 1049.500000 302.350000 ;
      RECT 957.500000 301.650000 999.500000 302.350000 ;
      RECT 907.500000 301.650000 949.500000 302.350000 ;
      RECT 857.500000 301.650000 899.500000 302.350000 ;
      RECT 807.500000 301.650000 849.500000 302.350000 ;
      RECT 757.500000 301.650000 799.500000 302.350000 ;
      RECT 707.500000 301.650000 749.500000 302.350000 ;
      RECT 657.500000 301.650000 699.500000 302.350000 ;
      RECT 607.500000 301.650000 649.500000 302.350000 ;
      RECT 557.500000 301.650000 599.500000 302.350000 ;
      RECT 507.500000 301.650000 549.500000 302.350000 ;
      RECT 407.500000 301.650000 458.500000 302.350000 ;
      RECT 357.500000 301.650000 399.500000 302.350000 ;
      RECT 307.500000 301.650000 349.500000 302.350000 ;
      RECT 257.500000 301.650000 299.500000 302.350000 ;
      RECT 207.500000 301.650000 249.500000 302.350000 ;
      RECT 157.500000 301.650000 199.500000 302.350000 ;
      RECT 107.500000 301.650000 149.500000 302.350000 ;
      RECT 57.500000 301.650000 99.500000 302.350000 ;
      RECT 15.500000 301.650000 49.500000 302.350000 ;
      RECT 1183.500000 300.350000 1186.000000 303.650000 ;
      RECT 1169.500000 300.350000 1170.500000 301.650000 ;
      RECT 1116.500000 300.350000 1149.500000 301.650000 ;
      RECT 1107.500000 300.350000 1108.500000 301.650000 ;
      RECT 1066.500000 300.350000 1099.500000 301.650000 ;
      RECT 1057.500000 300.350000 1058.500000 301.650000 ;
      RECT 1016.500000 300.350000 1049.500000 301.650000 ;
      RECT 1007.500000 300.350000 1008.500000 301.650000 ;
      RECT 966.500000 300.350000 999.500000 301.650000 ;
      RECT 957.500000 300.350000 958.500000 301.650000 ;
      RECT 916.500000 300.350000 949.500000 301.650000 ;
      RECT 907.500000 300.350000 908.500000 301.650000 ;
      RECT 866.500000 300.350000 899.500000 301.650000 ;
      RECT 857.500000 300.350000 858.500000 301.650000 ;
      RECT 816.500000 300.350000 849.500000 301.650000 ;
      RECT 807.500000 300.350000 808.500000 301.650000 ;
      RECT 766.500000 300.350000 799.500000 301.650000 ;
      RECT 757.500000 300.350000 758.500000 301.650000 ;
      RECT 716.500000 300.350000 749.500000 301.650000 ;
      RECT 707.500000 300.350000 708.500000 301.650000 ;
      RECT 666.500000 300.350000 699.500000 301.650000 ;
      RECT 657.500000 300.350000 658.500000 301.650000 ;
      RECT 616.500000 300.350000 649.500000 301.650000 ;
      RECT 607.500000 300.350000 608.500000 301.650000 ;
      RECT 566.500000 300.350000 599.500000 301.650000 ;
      RECT 557.500000 300.350000 558.500000 301.650000 ;
      RECT 516.500000 300.350000 549.500000 301.650000 ;
      RECT 507.500000 300.350000 508.500000 301.650000 ;
      RECT 466.500000 300.350000 499.500000 303.650000 ;
      RECT 407.500000 300.350000 408.500000 301.650000 ;
      RECT 366.500000 300.350000 399.500000 301.650000 ;
      RECT 357.500000 300.350000 358.500000 301.650000 ;
      RECT 316.500000 300.350000 349.500000 301.650000 ;
      RECT 307.500000 300.350000 308.500000 301.650000 ;
      RECT 266.500000 300.350000 299.500000 301.650000 ;
      RECT 257.500000 300.350000 258.500000 301.650000 ;
      RECT 216.500000 300.350000 249.500000 301.650000 ;
      RECT 207.500000 300.350000 208.500000 301.650000 ;
      RECT 166.500000 300.350000 199.500000 301.650000 ;
      RECT 157.500000 300.350000 158.500000 301.650000 ;
      RECT 116.500000 300.350000 149.500000 301.650000 ;
      RECT 107.500000 300.350000 108.500000 301.650000 ;
      RECT 66.500000 300.350000 99.500000 301.650000 ;
      RECT 57.500000 300.350000 58.500000 301.650000 ;
      RECT 29.500000 300.350000 49.500000 301.650000 ;
      RECT 15.500000 300.350000 16.500000 301.650000 ;
      RECT 0.000000 300.350000 2.500000 303.650000 ;
      RECT 466.500000 299.730000 508.500000 300.350000 ;
      RECT 416.500000 299.730000 458.500000 301.650000 ;
      RECT 1169.500000 299.650000 1186.000000 300.350000 ;
      RECT 1116.500000 299.650000 1156.500000 300.350000 ;
      RECT 1066.500000 299.650000 1108.500000 300.350000 ;
      RECT 1016.500000 299.650000 1058.500000 300.350000 ;
      RECT 966.500000 299.650000 1008.500000 300.350000 ;
      RECT 916.500000 299.650000 958.500000 300.350000 ;
      RECT 866.500000 299.650000 908.500000 300.350000 ;
      RECT 816.500000 299.650000 858.500000 300.350000 ;
      RECT 766.500000 299.650000 808.500000 300.350000 ;
      RECT 716.500000 299.650000 758.500000 300.350000 ;
      RECT 666.500000 299.650000 708.500000 300.350000 ;
      RECT 616.500000 299.650000 658.500000 300.350000 ;
      RECT 566.500000 299.650000 608.500000 300.350000 ;
      RECT 516.500000 299.650000 558.500000 300.350000 ;
      RECT 416.500000 299.650000 508.500000 299.730000 ;
      RECT 366.500000 299.650000 408.500000 300.350000 ;
      RECT 316.500000 299.650000 358.500000 300.350000 ;
      RECT 266.500000 299.650000 308.500000 300.350000 ;
      RECT 216.500000 299.650000 258.500000 300.350000 ;
      RECT 166.500000 299.650000 208.500000 300.350000 ;
      RECT 116.500000 299.650000 158.500000 300.350000 ;
      RECT 66.500000 299.650000 108.500000 300.350000 ;
      RECT 29.500000 299.650000 58.500000 300.350000 ;
      RECT 0.000000 299.650000 16.500000 300.350000 ;
      RECT 1169.500000 298.350000 1170.500000 299.650000 ;
      RECT 1116.500000 298.350000 1149.500000 299.650000 ;
      RECT 1107.500000 298.350000 1108.500000 299.650000 ;
      RECT 1066.500000 298.350000 1099.500000 299.650000 ;
      RECT 1057.500000 298.350000 1058.500000 299.650000 ;
      RECT 1016.500000 298.350000 1049.500000 299.650000 ;
      RECT 1007.500000 298.350000 1008.500000 299.650000 ;
      RECT 966.500000 298.350000 999.500000 299.650000 ;
      RECT 957.500000 298.350000 958.500000 299.650000 ;
      RECT 916.500000 298.350000 949.500000 299.650000 ;
      RECT 907.500000 298.350000 908.500000 299.650000 ;
      RECT 866.500000 298.350000 899.500000 299.650000 ;
      RECT 857.500000 298.350000 858.500000 299.650000 ;
      RECT 816.500000 298.350000 849.500000 299.650000 ;
      RECT 807.500000 298.350000 808.500000 299.650000 ;
      RECT 766.500000 298.350000 799.500000 299.650000 ;
      RECT 757.500000 298.350000 758.500000 299.650000 ;
      RECT 716.500000 298.350000 749.500000 299.650000 ;
      RECT 707.500000 298.350000 708.500000 299.650000 ;
      RECT 666.500000 298.350000 699.500000 299.650000 ;
      RECT 657.500000 298.350000 658.500000 299.650000 ;
      RECT 616.500000 298.350000 649.500000 299.650000 ;
      RECT 607.500000 298.350000 608.500000 299.650000 ;
      RECT 566.500000 298.350000 599.500000 299.650000 ;
      RECT 557.500000 298.350000 558.500000 299.650000 ;
      RECT 516.500000 298.350000 549.500000 299.650000 ;
      RECT 507.500000 298.350000 508.500000 299.650000 ;
      RECT 416.500000 298.350000 449.500000 299.650000 ;
      RECT 407.500000 298.350000 408.500000 299.650000 ;
      RECT 366.500000 298.350000 399.500000 299.650000 ;
      RECT 357.500000 298.350000 358.500000 299.650000 ;
      RECT 316.500000 298.350000 349.500000 299.650000 ;
      RECT 307.500000 298.350000 308.500000 299.650000 ;
      RECT 266.500000 298.350000 299.500000 299.650000 ;
      RECT 257.500000 298.350000 258.500000 299.650000 ;
      RECT 216.500000 298.350000 249.500000 299.650000 ;
      RECT 207.500000 298.350000 208.500000 299.650000 ;
      RECT 166.500000 298.350000 199.500000 299.650000 ;
      RECT 157.500000 298.350000 158.500000 299.650000 ;
      RECT 116.500000 298.350000 149.500000 299.650000 ;
      RECT 107.500000 298.350000 108.500000 299.650000 ;
      RECT 66.500000 298.350000 99.500000 299.650000 ;
      RECT 57.500000 298.350000 58.500000 299.650000 ;
      RECT 29.500000 298.350000 49.500000 299.650000 ;
      RECT 15.500000 298.350000 16.500000 299.650000 ;
      RECT 1157.500000 297.650000 1170.500000 298.350000 ;
      RECT 1107.500000 297.650000 1149.500000 298.350000 ;
      RECT 1057.500000 297.650000 1099.500000 298.350000 ;
      RECT 1007.500000 297.650000 1049.500000 298.350000 ;
      RECT 957.500000 297.650000 999.500000 298.350000 ;
      RECT 907.500000 297.650000 949.500000 298.350000 ;
      RECT 857.500000 297.650000 899.500000 298.350000 ;
      RECT 807.500000 297.650000 849.500000 298.350000 ;
      RECT 757.500000 297.650000 799.500000 298.350000 ;
      RECT 707.500000 297.650000 749.500000 298.350000 ;
      RECT 657.500000 297.650000 699.500000 298.350000 ;
      RECT 607.500000 297.650000 649.500000 298.350000 ;
      RECT 557.500000 297.650000 599.500000 298.350000 ;
      RECT 507.500000 297.650000 549.500000 298.350000 ;
      RECT 457.500000 297.650000 499.500000 299.650000 ;
      RECT 407.500000 297.650000 449.500000 298.350000 ;
      RECT 357.500000 297.650000 399.500000 298.350000 ;
      RECT 307.500000 297.650000 349.500000 298.350000 ;
      RECT 257.500000 297.650000 299.500000 298.350000 ;
      RECT 207.500000 297.650000 249.500000 298.350000 ;
      RECT 157.500000 297.650000 199.500000 298.350000 ;
      RECT 107.500000 297.650000 149.500000 298.350000 ;
      RECT 57.500000 297.650000 99.500000 298.350000 ;
      RECT 15.500000 297.650000 49.500000 298.350000 ;
      RECT 1183.500000 296.350000 1186.000000 299.650000 ;
      RECT 1169.500000 296.350000 1170.500000 297.650000 ;
      RECT 1116.500000 296.350000 1149.500000 297.650000 ;
      RECT 1107.500000 296.350000 1108.500000 297.650000 ;
      RECT 1066.500000 296.350000 1099.500000 297.650000 ;
      RECT 1057.500000 296.350000 1058.500000 297.650000 ;
      RECT 1016.500000 296.350000 1049.500000 297.650000 ;
      RECT 1007.500000 296.350000 1008.500000 297.650000 ;
      RECT 966.500000 296.350000 999.500000 297.650000 ;
      RECT 957.500000 296.350000 958.500000 297.650000 ;
      RECT 916.500000 296.350000 949.500000 297.650000 ;
      RECT 907.500000 296.350000 908.500000 297.650000 ;
      RECT 866.500000 296.350000 899.500000 297.650000 ;
      RECT 857.500000 296.350000 858.500000 297.650000 ;
      RECT 816.500000 296.350000 849.500000 297.650000 ;
      RECT 807.500000 296.350000 808.500000 297.650000 ;
      RECT 766.500000 296.350000 799.500000 297.650000 ;
      RECT 757.500000 296.350000 758.500000 297.650000 ;
      RECT 716.500000 296.350000 749.500000 297.650000 ;
      RECT 707.500000 296.350000 708.500000 297.650000 ;
      RECT 666.500000 296.350000 699.500000 297.650000 ;
      RECT 657.500000 296.350000 658.500000 297.650000 ;
      RECT 616.500000 296.350000 649.500000 297.650000 ;
      RECT 607.500000 296.350000 608.500000 297.650000 ;
      RECT 566.500000 296.350000 599.500000 297.650000 ;
      RECT 557.500000 296.350000 558.500000 297.650000 ;
      RECT 516.500000 296.350000 549.500000 297.650000 ;
      RECT 507.500000 296.350000 508.500000 297.650000 ;
      RECT 466.500000 296.350000 499.500000 297.650000 ;
      RECT 457.500000 296.350000 458.500000 297.650000 ;
      RECT 416.500000 296.350000 449.500000 297.650000 ;
      RECT 407.500000 296.350000 408.500000 297.650000 ;
      RECT 366.500000 296.350000 399.500000 297.650000 ;
      RECT 357.500000 296.350000 358.500000 297.650000 ;
      RECT 316.500000 296.350000 349.500000 297.650000 ;
      RECT 307.500000 296.350000 308.500000 297.650000 ;
      RECT 266.500000 296.350000 299.500000 297.650000 ;
      RECT 257.500000 296.350000 258.500000 297.650000 ;
      RECT 216.500000 296.350000 249.500000 297.650000 ;
      RECT 207.500000 296.350000 208.500000 297.650000 ;
      RECT 166.500000 296.350000 199.500000 297.650000 ;
      RECT 157.500000 296.350000 158.500000 297.650000 ;
      RECT 116.500000 296.350000 149.500000 297.650000 ;
      RECT 107.500000 296.350000 108.500000 297.650000 ;
      RECT 66.500000 296.350000 99.500000 297.650000 ;
      RECT 57.500000 296.350000 58.500000 297.650000 ;
      RECT 29.500000 296.350000 49.500000 297.650000 ;
      RECT 15.500000 296.350000 16.500000 297.650000 ;
      RECT 0.000000 296.350000 2.500000 299.650000 ;
      RECT 1169.500000 295.650000 1186.000000 296.350000 ;
      RECT 1116.500000 295.650000 1156.500000 296.350000 ;
      RECT 1066.500000 295.650000 1108.500000 296.350000 ;
      RECT 1016.500000 295.650000 1058.500000 296.350000 ;
      RECT 966.500000 295.650000 1008.500000 296.350000 ;
      RECT 916.500000 295.650000 958.500000 296.350000 ;
      RECT 866.500000 295.650000 908.500000 296.350000 ;
      RECT 816.500000 295.650000 858.500000 296.350000 ;
      RECT 766.500000 295.650000 808.500000 296.350000 ;
      RECT 716.500000 295.650000 758.500000 296.350000 ;
      RECT 666.500000 295.650000 708.500000 296.350000 ;
      RECT 616.500000 295.650000 658.500000 296.350000 ;
      RECT 566.500000 295.650000 608.500000 296.350000 ;
      RECT 516.500000 295.650000 558.500000 296.350000 ;
      RECT 466.500000 295.650000 508.500000 296.350000 ;
      RECT 416.500000 295.650000 458.500000 296.350000 ;
      RECT 366.500000 295.650000 408.500000 296.350000 ;
      RECT 316.500000 295.650000 358.500000 296.350000 ;
      RECT 266.500000 295.650000 308.500000 296.350000 ;
      RECT 216.500000 295.650000 258.500000 296.350000 ;
      RECT 166.500000 295.650000 208.500000 296.350000 ;
      RECT 116.500000 295.650000 158.500000 296.350000 ;
      RECT 66.500000 295.650000 108.500000 296.350000 ;
      RECT 29.500000 295.650000 58.500000 296.350000 ;
      RECT 0.000000 295.650000 16.500000 296.350000 ;
      RECT 1169.500000 294.350000 1170.500000 295.650000 ;
      RECT 1116.500000 294.350000 1149.500000 295.650000 ;
      RECT 1107.500000 294.350000 1108.500000 295.650000 ;
      RECT 1066.500000 294.350000 1099.500000 295.650000 ;
      RECT 1057.500000 294.350000 1058.500000 295.650000 ;
      RECT 1016.500000 294.350000 1049.500000 295.650000 ;
      RECT 1007.500000 294.350000 1008.500000 295.650000 ;
      RECT 966.500000 294.350000 999.500000 295.650000 ;
      RECT 957.500000 294.350000 958.500000 295.650000 ;
      RECT 916.500000 294.350000 949.500000 295.650000 ;
      RECT 907.500000 294.350000 908.500000 295.650000 ;
      RECT 866.500000 294.350000 899.500000 295.650000 ;
      RECT 857.500000 294.350000 858.500000 295.650000 ;
      RECT 816.500000 294.350000 849.500000 295.650000 ;
      RECT 807.500000 294.350000 808.500000 295.650000 ;
      RECT 766.500000 294.350000 799.500000 295.650000 ;
      RECT 757.500000 294.350000 758.500000 295.650000 ;
      RECT 716.500000 294.350000 749.500000 295.650000 ;
      RECT 707.500000 294.350000 708.500000 295.650000 ;
      RECT 666.500000 294.350000 699.500000 295.650000 ;
      RECT 657.500000 294.350000 658.500000 295.650000 ;
      RECT 616.500000 294.350000 649.500000 295.650000 ;
      RECT 607.500000 294.350000 608.500000 295.650000 ;
      RECT 566.500000 294.350000 599.500000 295.650000 ;
      RECT 557.500000 294.350000 558.500000 295.650000 ;
      RECT 516.500000 294.350000 549.500000 295.650000 ;
      RECT 507.500000 294.350000 508.500000 295.650000 ;
      RECT 466.500000 294.350000 499.500000 295.650000 ;
      RECT 457.500000 294.350000 458.500000 295.650000 ;
      RECT 416.500000 294.350000 449.500000 295.650000 ;
      RECT 407.500000 294.350000 408.500000 295.650000 ;
      RECT 366.500000 294.350000 399.500000 295.650000 ;
      RECT 357.500000 294.350000 358.500000 295.650000 ;
      RECT 316.500000 294.350000 349.500000 295.650000 ;
      RECT 307.500000 294.350000 308.500000 295.650000 ;
      RECT 266.500000 294.350000 299.500000 295.650000 ;
      RECT 257.500000 294.350000 258.500000 295.650000 ;
      RECT 216.500000 294.350000 249.500000 295.650000 ;
      RECT 207.500000 294.350000 208.500000 295.650000 ;
      RECT 166.500000 294.350000 199.500000 295.650000 ;
      RECT 157.500000 294.350000 158.500000 295.650000 ;
      RECT 116.500000 294.350000 149.500000 295.650000 ;
      RECT 107.500000 294.350000 108.500000 295.650000 ;
      RECT 66.500000 294.350000 99.500000 295.650000 ;
      RECT 57.500000 294.350000 58.500000 295.650000 ;
      RECT 29.500000 294.350000 49.500000 295.650000 ;
      RECT 15.500000 294.350000 16.500000 295.650000 ;
      RECT 1157.500000 293.650000 1170.500000 294.350000 ;
      RECT 1107.500000 293.650000 1149.500000 294.350000 ;
      RECT 1057.500000 293.650000 1099.500000 294.350000 ;
      RECT 1007.500000 293.650000 1049.500000 294.350000 ;
      RECT 957.500000 293.650000 999.500000 294.350000 ;
      RECT 907.500000 293.650000 949.500000 294.350000 ;
      RECT 857.500000 293.650000 899.500000 294.350000 ;
      RECT 807.500000 293.650000 849.500000 294.350000 ;
      RECT 757.500000 293.650000 799.500000 294.350000 ;
      RECT 707.500000 293.650000 749.500000 294.350000 ;
      RECT 657.500000 293.650000 699.500000 294.350000 ;
      RECT 607.500000 293.650000 649.500000 294.350000 ;
      RECT 557.500000 293.650000 599.500000 294.350000 ;
      RECT 507.500000 293.650000 549.500000 294.350000 ;
      RECT 457.500000 293.650000 499.500000 294.350000 ;
      RECT 407.500000 293.650000 449.500000 294.350000 ;
      RECT 357.500000 293.650000 399.500000 294.350000 ;
      RECT 307.500000 293.650000 349.500000 294.350000 ;
      RECT 257.500000 293.650000 299.500000 294.350000 ;
      RECT 207.500000 293.650000 249.500000 294.350000 ;
      RECT 157.500000 293.650000 199.500000 294.350000 ;
      RECT 107.500000 293.650000 149.500000 294.350000 ;
      RECT 57.500000 293.650000 99.500000 294.350000 ;
      RECT 15.500000 293.650000 49.500000 294.350000 ;
      RECT 1183.500000 292.350000 1186.000000 295.650000 ;
      RECT 1169.500000 292.350000 1170.500000 293.650000 ;
      RECT 1116.500000 292.350000 1149.500000 293.650000 ;
      RECT 1107.500000 292.350000 1108.500000 293.650000 ;
      RECT 1066.500000 292.350000 1099.500000 293.650000 ;
      RECT 1057.500000 292.350000 1058.500000 293.650000 ;
      RECT 1016.500000 292.350000 1049.500000 293.650000 ;
      RECT 1007.500000 292.350000 1008.500000 293.650000 ;
      RECT 966.500000 292.350000 999.500000 293.650000 ;
      RECT 957.500000 292.350000 958.500000 293.650000 ;
      RECT 916.500000 292.350000 949.500000 293.650000 ;
      RECT 907.500000 292.350000 908.500000 293.650000 ;
      RECT 866.500000 292.350000 899.500000 293.650000 ;
      RECT 857.500000 292.350000 858.500000 293.650000 ;
      RECT 816.500000 292.350000 849.500000 293.650000 ;
      RECT 807.500000 292.350000 808.500000 293.650000 ;
      RECT 766.500000 292.350000 799.500000 293.650000 ;
      RECT 757.500000 292.350000 758.500000 293.650000 ;
      RECT 716.500000 292.350000 749.500000 293.650000 ;
      RECT 707.500000 292.350000 708.500000 293.650000 ;
      RECT 666.500000 292.350000 699.500000 293.650000 ;
      RECT 657.500000 292.350000 658.500000 293.650000 ;
      RECT 616.500000 292.350000 649.500000 293.650000 ;
      RECT 607.500000 292.350000 608.500000 293.650000 ;
      RECT 566.500000 292.350000 599.500000 293.650000 ;
      RECT 557.500000 292.350000 558.500000 293.650000 ;
      RECT 516.500000 292.350000 549.500000 293.650000 ;
      RECT 507.500000 292.350000 508.500000 293.650000 ;
      RECT 466.500000 292.350000 499.500000 293.650000 ;
      RECT 457.500000 292.350000 458.500000 293.650000 ;
      RECT 416.500000 292.350000 449.500000 293.650000 ;
      RECT 407.500000 292.350000 408.500000 293.650000 ;
      RECT 366.500000 292.350000 399.500000 293.650000 ;
      RECT 357.500000 292.350000 358.500000 293.650000 ;
      RECT 316.500000 292.350000 349.500000 293.650000 ;
      RECT 307.500000 292.350000 308.500000 293.650000 ;
      RECT 266.500000 292.350000 299.500000 293.650000 ;
      RECT 257.500000 292.350000 258.500000 293.650000 ;
      RECT 216.500000 292.350000 249.500000 293.650000 ;
      RECT 207.500000 292.350000 208.500000 293.650000 ;
      RECT 166.500000 292.350000 199.500000 293.650000 ;
      RECT 157.500000 292.350000 158.500000 293.650000 ;
      RECT 116.500000 292.350000 149.500000 293.650000 ;
      RECT 107.500000 292.350000 108.500000 293.650000 ;
      RECT 66.500000 292.350000 99.500000 293.650000 ;
      RECT 57.500000 292.350000 58.500000 293.650000 ;
      RECT 29.500000 292.350000 49.500000 293.650000 ;
      RECT 15.500000 292.350000 16.500000 293.650000 ;
      RECT 0.000000 292.350000 2.500000 295.650000 ;
      RECT 1169.500000 291.650000 1186.000000 292.350000 ;
      RECT 1116.500000 291.650000 1156.500000 292.350000 ;
      RECT 1066.500000 291.650000 1108.500000 292.350000 ;
      RECT 1016.500000 291.650000 1058.500000 292.350000 ;
      RECT 966.500000 291.650000 1008.500000 292.350000 ;
      RECT 916.500000 291.650000 958.500000 292.350000 ;
      RECT 866.500000 291.650000 908.500000 292.350000 ;
      RECT 816.500000 291.650000 858.500000 292.350000 ;
      RECT 766.500000 291.650000 808.500000 292.350000 ;
      RECT 716.500000 291.650000 758.500000 292.350000 ;
      RECT 666.500000 291.650000 708.500000 292.350000 ;
      RECT 616.500000 291.650000 658.500000 292.350000 ;
      RECT 566.500000 291.650000 608.500000 292.350000 ;
      RECT 516.500000 291.650000 558.500000 292.350000 ;
      RECT 466.500000 291.650000 508.500000 292.350000 ;
      RECT 416.500000 291.650000 458.500000 292.350000 ;
      RECT 366.500000 291.650000 408.500000 292.350000 ;
      RECT 316.500000 291.650000 358.500000 292.350000 ;
      RECT 266.500000 291.650000 308.500000 292.350000 ;
      RECT 216.500000 291.650000 258.500000 292.350000 ;
      RECT 166.500000 291.650000 208.500000 292.350000 ;
      RECT 116.500000 291.650000 158.500000 292.350000 ;
      RECT 66.500000 291.650000 108.500000 292.350000 ;
      RECT 29.500000 291.650000 58.500000 292.350000 ;
      RECT 0.000000 291.650000 16.500000 292.350000 ;
      RECT 1169.500000 290.350000 1170.500000 291.650000 ;
      RECT 1116.500000 290.350000 1149.500000 291.650000 ;
      RECT 1107.500000 290.350000 1108.500000 291.650000 ;
      RECT 1066.500000 290.350000 1099.500000 291.650000 ;
      RECT 1057.500000 290.350000 1058.500000 291.650000 ;
      RECT 1016.500000 290.350000 1049.500000 291.650000 ;
      RECT 1007.500000 290.350000 1008.500000 291.650000 ;
      RECT 966.500000 290.350000 999.500000 291.650000 ;
      RECT 957.500000 290.350000 958.500000 291.650000 ;
      RECT 916.500000 290.350000 949.500000 291.650000 ;
      RECT 907.500000 290.350000 908.500000 291.650000 ;
      RECT 866.500000 290.350000 899.500000 291.650000 ;
      RECT 857.500000 290.350000 858.500000 291.650000 ;
      RECT 816.500000 290.350000 849.500000 291.650000 ;
      RECT 807.500000 290.350000 808.500000 291.650000 ;
      RECT 766.500000 290.350000 799.500000 291.650000 ;
      RECT 757.500000 290.350000 758.500000 291.650000 ;
      RECT 716.500000 290.350000 749.500000 291.650000 ;
      RECT 707.500000 290.350000 708.500000 291.650000 ;
      RECT 666.500000 290.350000 699.500000 291.650000 ;
      RECT 657.500000 290.350000 658.500000 291.650000 ;
      RECT 616.500000 290.350000 649.500000 291.650000 ;
      RECT 607.500000 290.350000 608.500000 291.650000 ;
      RECT 566.500000 290.350000 599.500000 291.650000 ;
      RECT 557.500000 290.350000 558.500000 291.650000 ;
      RECT 516.500000 290.350000 549.500000 291.650000 ;
      RECT 507.500000 290.350000 508.500000 291.650000 ;
      RECT 466.500000 290.350000 499.500000 291.650000 ;
      RECT 457.500000 290.350000 458.500000 291.650000 ;
      RECT 416.500000 290.350000 449.500000 291.650000 ;
      RECT 407.500000 290.350000 408.500000 291.650000 ;
      RECT 366.500000 290.350000 399.500000 291.650000 ;
      RECT 357.500000 290.350000 358.500000 291.650000 ;
      RECT 316.500000 290.350000 349.500000 291.650000 ;
      RECT 307.500000 290.350000 308.500000 291.650000 ;
      RECT 266.500000 290.350000 299.500000 291.650000 ;
      RECT 257.500000 290.350000 258.500000 291.650000 ;
      RECT 216.500000 290.350000 249.500000 291.650000 ;
      RECT 207.500000 290.350000 208.500000 291.650000 ;
      RECT 166.500000 290.350000 199.500000 291.650000 ;
      RECT 157.500000 290.350000 158.500000 291.650000 ;
      RECT 116.500000 290.350000 149.500000 291.650000 ;
      RECT 107.500000 290.350000 108.500000 291.650000 ;
      RECT 66.500000 290.350000 99.500000 291.650000 ;
      RECT 57.500000 290.350000 58.500000 291.650000 ;
      RECT 29.500000 290.350000 49.500000 291.650000 ;
      RECT 15.500000 290.350000 16.500000 291.650000 ;
      RECT 1157.500000 289.650000 1170.500000 290.350000 ;
      RECT 1107.500000 289.650000 1149.500000 290.350000 ;
      RECT 1057.500000 289.650000 1099.500000 290.350000 ;
      RECT 1007.500000 289.650000 1049.500000 290.350000 ;
      RECT 957.500000 289.650000 999.500000 290.350000 ;
      RECT 907.500000 289.650000 949.500000 290.350000 ;
      RECT 857.500000 289.650000 899.500000 290.350000 ;
      RECT 807.500000 289.650000 849.500000 290.350000 ;
      RECT 757.500000 289.650000 799.500000 290.350000 ;
      RECT 707.500000 289.650000 749.500000 290.350000 ;
      RECT 657.500000 289.650000 699.500000 290.350000 ;
      RECT 607.500000 289.650000 649.500000 290.350000 ;
      RECT 557.500000 289.650000 599.500000 290.350000 ;
      RECT 507.500000 289.650000 549.500000 290.350000 ;
      RECT 457.500000 289.650000 499.500000 290.350000 ;
      RECT 407.500000 289.650000 449.500000 290.350000 ;
      RECT 357.500000 289.650000 399.500000 290.350000 ;
      RECT 307.500000 289.650000 349.500000 290.350000 ;
      RECT 257.500000 289.650000 299.500000 290.350000 ;
      RECT 207.500000 289.650000 249.500000 290.350000 ;
      RECT 157.500000 289.650000 199.500000 290.350000 ;
      RECT 107.500000 289.650000 149.500000 290.350000 ;
      RECT 57.500000 289.650000 99.500000 290.350000 ;
      RECT 15.500000 289.650000 49.500000 290.350000 ;
      RECT 1183.500000 288.350000 1186.000000 291.650000 ;
      RECT 1169.500000 288.350000 1170.500000 289.650000 ;
      RECT 1116.500000 288.350000 1149.500000 289.650000 ;
      RECT 1107.500000 288.350000 1108.500000 289.650000 ;
      RECT 1066.500000 288.350000 1099.500000 289.650000 ;
      RECT 1057.500000 288.350000 1058.500000 289.650000 ;
      RECT 1016.500000 288.350000 1049.500000 289.650000 ;
      RECT 1007.500000 288.350000 1008.500000 289.650000 ;
      RECT 966.500000 288.350000 999.500000 289.650000 ;
      RECT 957.500000 288.350000 958.500000 289.650000 ;
      RECT 916.500000 288.350000 949.500000 289.650000 ;
      RECT 907.500000 288.350000 908.500000 289.650000 ;
      RECT 866.500000 288.350000 899.500000 289.650000 ;
      RECT 857.500000 288.350000 858.500000 289.650000 ;
      RECT 816.500000 288.350000 849.500000 289.650000 ;
      RECT 807.500000 288.350000 808.500000 289.650000 ;
      RECT 766.500000 288.350000 799.500000 289.650000 ;
      RECT 757.500000 288.350000 758.500000 289.650000 ;
      RECT 716.500000 288.350000 749.500000 289.650000 ;
      RECT 707.500000 288.350000 708.500000 289.650000 ;
      RECT 666.500000 288.350000 699.500000 289.650000 ;
      RECT 657.500000 288.350000 658.500000 289.650000 ;
      RECT 616.500000 288.350000 649.500000 289.650000 ;
      RECT 607.500000 288.350000 608.500000 289.650000 ;
      RECT 566.500000 288.350000 599.500000 289.650000 ;
      RECT 557.500000 288.350000 558.500000 289.650000 ;
      RECT 516.500000 288.350000 549.500000 289.650000 ;
      RECT 507.500000 288.350000 508.500000 289.650000 ;
      RECT 466.500000 288.350000 499.500000 289.650000 ;
      RECT 457.500000 288.350000 458.500000 289.650000 ;
      RECT 416.500000 288.350000 449.500000 289.650000 ;
      RECT 407.500000 288.350000 408.500000 289.650000 ;
      RECT 366.500000 288.350000 399.500000 289.650000 ;
      RECT 357.500000 288.350000 358.500000 289.650000 ;
      RECT 316.500000 288.350000 349.500000 289.650000 ;
      RECT 307.500000 288.350000 308.500000 289.650000 ;
      RECT 266.500000 288.350000 299.500000 289.650000 ;
      RECT 257.500000 288.350000 258.500000 289.650000 ;
      RECT 216.500000 288.350000 249.500000 289.650000 ;
      RECT 207.500000 288.350000 208.500000 289.650000 ;
      RECT 166.500000 288.350000 199.500000 289.650000 ;
      RECT 157.500000 288.350000 158.500000 289.650000 ;
      RECT 116.500000 288.350000 149.500000 289.650000 ;
      RECT 107.500000 288.350000 108.500000 289.650000 ;
      RECT 66.500000 288.350000 99.500000 289.650000 ;
      RECT 57.500000 288.350000 58.500000 289.650000 ;
      RECT 29.500000 288.350000 49.500000 289.650000 ;
      RECT 15.500000 288.350000 16.500000 289.650000 ;
      RECT 0.000000 288.350000 2.500000 291.650000 ;
      RECT 1169.500000 287.650000 1186.000000 288.350000 ;
      RECT 1116.500000 287.650000 1156.500000 288.350000 ;
      RECT 1066.500000 287.650000 1108.500000 288.350000 ;
      RECT 1016.500000 287.650000 1058.500000 288.350000 ;
      RECT 966.500000 287.650000 1008.500000 288.350000 ;
      RECT 916.500000 287.650000 958.500000 288.350000 ;
      RECT 866.500000 287.650000 908.500000 288.350000 ;
      RECT 816.500000 287.650000 858.500000 288.350000 ;
      RECT 766.500000 287.650000 808.500000 288.350000 ;
      RECT 716.500000 287.650000 758.500000 288.350000 ;
      RECT 666.500000 287.650000 708.500000 288.350000 ;
      RECT 616.500000 287.650000 658.500000 288.350000 ;
      RECT 566.500000 287.650000 608.500000 288.350000 ;
      RECT 516.500000 287.650000 558.500000 288.350000 ;
      RECT 466.500000 287.650000 508.500000 288.350000 ;
      RECT 416.500000 287.650000 458.500000 288.350000 ;
      RECT 366.500000 287.650000 408.500000 288.350000 ;
      RECT 316.500000 287.650000 358.500000 288.350000 ;
      RECT 266.500000 287.650000 308.500000 288.350000 ;
      RECT 216.500000 287.650000 258.500000 288.350000 ;
      RECT 166.500000 287.650000 208.500000 288.350000 ;
      RECT 116.500000 287.650000 158.500000 288.350000 ;
      RECT 66.500000 287.650000 108.500000 288.350000 ;
      RECT 29.500000 287.650000 58.500000 288.350000 ;
      RECT 0.000000 287.650000 16.500000 288.350000 ;
      RECT 1169.500000 286.350000 1170.500000 287.650000 ;
      RECT 1116.500000 286.350000 1149.500000 287.650000 ;
      RECT 1107.500000 286.350000 1108.500000 287.650000 ;
      RECT 1066.500000 286.350000 1099.500000 287.650000 ;
      RECT 1057.500000 286.350000 1058.500000 287.650000 ;
      RECT 1016.500000 286.350000 1049.500000 287.650000 ;
      RECT 1007.500000 286.350000 1008.500000 287.650000 ;
      RECT 966.500000 286.350000 999.500000 287.650000 ;
      RECT 957.500000 286.350000 958.500000 287.650000 ;
      RECT 916.500000 286.350000 949.500000 287.650000 ;
      RECT 907.500000 286.350000 908.500000 287.650000 ;
      RECT 866.500000 286.350000 899.500000 287.650000 ;
      RECT 857.500000 286.350000 858.500000 287.650000 ;
      RECT 816.500000 286.350000 849.500000 287.650000 ;
      RECT 807.500000 286.350000 808.500000 287.650000 ;
      RECT 766.500000 286.350000 799.500000 287.650000 ;
      RECT 757.500000 286.350000 758.500000 287.650000 ;
      RECT 716.500000 286.350000 749.500000 287.650000 ;
      RECT 707.500000 286.350000 708.500000 287.650000 ;
      RECT 666.500000 286.350000 699.500000 287.650000 ;
      RECT 657.500000 286.350000 658.500000 287.650000 ;
      RECT 616.500000 286.350000 649.500000 287.650000 ;
      RECT 607.500000 286.350000 608.500000 287.650000 ;
      RECT 566.500000 286.350000 599.500000 287.650000 ;
      RECT 557.500000 286.350000 558.500000 287.650000 ;
      RECT 516.500000 286.350000 549.500000 287.650000 ;
      RECT 507.500000 286.350000 508.500000 287.650000 ;
      RECT 466.500000 286.350000 499.500000 287.650000 ;
      RECT 457.500000 286.350000 458.500000 287.650000 ;
      RECT 416.500000 286.350000 449.500000 287.650000 ;
      RECT 407.500000 286.350000 408.500000 287.650000 ;
      RECT 366.500000 286.350000 399.500000 287.650000 ;
      RECT 357.500000 286.350000 358.500000 287.650000 ;
      RECT 316.500000 286.350000 349.500000 287.650000 ;
      RECT 307.500000 286.350000 308.500000 287.650000 ;
      RECT 266.500000 286.350000 299.500000 287.650000 ;
      RECT 257.500000 286.350000 258.500000 287.650000 ;
      RECT 216.500000 286.350000 249.500000 287.650000 ;
      RECT 207.500000 286.350000 208.500000 287.650000 ;
      RECT 166.500000 286.350000 199.500000 287.650000 ;
      RECT 157.500000 286.350000 158.500000 287.650000 ;
      RECT 116.500000 286.350000 149.500000 287.650000 ;
      RECT 107.500000 286.350000 108.500000 287.650000 ;
      RECT 66.500000 286.350000 99.500000 287.650000 ;
      RECT 57.500000 286.350000 58.500000 287.650000 ;
      RECT 29.500000 286.350000 49.500000 287.650000 ;
      RECT 15.500000 286.350000 16.500000 287.650000 ;
      RECT 1157.500000 285.650000 1170.500000 286.350000 ;
      RECT 1107.500000 285.650000 1149.500000 286.350000 ;
      RECT 1057.500000 285.650000 1099.500000 286.350000 ;
      RECT 1007.500000 285.650000 1049.500000 286.350000 ;
      RECT 957.500000 285.650000 999.500000 286.350000 ;
      RECT 907.500000 285.650000 949.500000 286.350000 ;
      RECT 857.500000 285.650000 899.500000 286.350000 ;
      RECT 807.500000 285.650000 849.500000 286.350000 ;
      RECT 757.500000 285.650000 799.500000 286.350000 ;
      RECT 707.500000 285.650000 749.500000 286.350000 ;
      RECT 657.500000 285.650000 699.500000 286.350000 ;
      RECT 607.500000 285.650000 649.500000 286.350000 ;
      RECT 557.500000 285.650000 599.500000 286.350000 ;
      RECT 507.500000 285.650000 549.500000 286.350000 ;
      RECT 457.500000 285.650000 499.500000 286.350000 ;
      RECT 407.500000 285.650000 449.500000 286.350000 ;
      RECT 357.500000 285.650000 399.500000 286.350000 ;
      RECT 307.500000 285.650000 349.500000 286.350000 ;
      RECT 257.500000 285.650000 299.500000 286.350000 ;
      RECT 207.500000 285.650000 249.500000 286.350000 ;
      RECT 157.500000 285.650000 199.500000 286.350000 ;
      RECT 107.500000 285.650000 149.500000 286.350000 ;
      RECT 57.500000 285.650000 99.500000 286.350000 ;
      RECT 15.500000 285.650000 49.500000 286.350000 ;
      RECT 1183.500000 284.350000 1186.000000 287.650000 ;
      RECT 1169.500000 284.350000 1170.500000 285.650000 ;
      RECT 1116.500000 284.350000 1149.500000 285.650000 ;
      RECT 1107.500000 284.350000 1108.500000 285.650000 ;
      RECT 1066.500000 284.350000 1099.500000 285.650000 ;
      RECT 1057.500000 284.350000 1058.500000 285.650000 ;
      RECT 1016.500000 284.350000 1049.500000 285.650000 ;
      RECT 1007.500000 284.350000 1008.500000 285.650000 ;
      RECT 966.500000 284.350000 999.500000 285.650000 ;
      RECT 957.500000 284.350000 958.500000 285.650000 ;
      RECT 916.500000 284.350000 949.500000 285.650000 ;
      RECT 907.500000 284.350000 908.500000 285.650000 ;
      RECT 866.500000 284.350000 899.500000 285.650000 ;
      RECT 857.500000 284.350000 858.500000 285.650000 ;
      RECT 816.500000 284.350000 849.500000 285.650000 ;
      RECT 807.500000 284.350000 808.500000 285.650000 ;
      RECT 766.500000 284.350000 799.500000 285.650000 ;
      RECT 757.500000 284.350000 758.500000 285.650000 ;
      RECT 716.500000 284.350000 749.500000 285.650000 ;
      RECT 707.500000 284.350000 708.500000 285.650000 ;
      RECT 666.500000 284.350000 699.500000 285.650000 ;
      RECT 657.500000 284.350000 658.500000 285.650000 ;
      RECT 616.500000 284.350000 649.500000 285.650000 ;
      RECT 607.500000 284.350000 608.500000 285.650000 ;
      RECT 566.500000 284.350000 599.500000 285.650000 ;
      RECT 557.500000 284.350000 558.500000 285.650000 ;
      RECT 516.500000 284.350000 549.500000 285.650000 ;
      RECT 507.500000 284.350000 508.500000 285.650000 ;
      RECT 466.500000 284.350000 499.500000 285.650000 ;
      RECT 457.500000 284.350000 458.500000 285.650000 ;
      RECT 416.500000 284.350000 449.500000 285.650000 ;
      RECT 407.500000 284.350000 408.500000 285.650000 ;
      RECT 366.500000 284.350000 399.500000 285.650000 ;
      RECT 357.500000 284.350000 358.500000 285.650000 ;
      RECT 316.500000 284.350000 349.500000 285.650000 ;
      RECT 307.500000 284.350000 308.500000 285.650000 ;
      RECT 266.500000 284.350000 299.500000 285.650000 ;
      RECT 257.500000 284.350000 258.500000 285.650000 ;
      RECT 216.500000 284.350000 249.500000 285.650000 ;
      RECT 207.500000 284.350000 208.500000 285.650000 ;
      RECT 166.500000 284.350000 199.500000 285.650000 ;
      RECT 157.500000 284.350000 158.500000 285.650000 ;
      RECT 116.500000 284.350000 149.500000 285.650000 ;
      RECT 107.500000 284.350000 108.500000 285.650000 ;
      RECT 66.500000 284.350000 99.500000 285.650000 ;
      RECT 57.500000 284.350000 58.500000 285.650000 ;
      RECT 29.500000 284.350000 49.500000 285.650000 ;
      RECT 15.500000 284.350000 16.500000 285.650000 ;
      RECT 0.000000 284.350000 2.500000 287.650000 ;
      RECT 1169.500000 283.650000 1186.000000 284.350000 ;
      RECT 1116.500000 283.650000 1156.500000 284.350000 ;
      RECT 1066.500000 283.650000 1108.500000 284.350000 ;
      RECT 1016.500000 283.650000 1058.500000 284.350000 ;
      RECT 966.500000 283.650000 1008.500000 284.350000 ;
      RECT 916.500000 283.650000 958.500000 284.350000 ;
      RECT 866.500000 283.650000 908.500000 284.350000 ;
      RECT 816.500000 283.650000 858.500000 284.350000 ;
      RECT 766.500000 283.650000 808.500000 284.350000 ;
      RECT 716.500000 283.650000 758.500000 284.350000 ;
      RECT 666.500000 283.650000 708.500000 284.350000 ;
      RECT 616.500000 283.650000 658.500000 284.350000 ;
      RECT 566.500000 283.650000 608.500000 284.350000 ;
      RECT 516.500000 283.650000 558.500000 284.350000 ;
      RECT 466.500000 283.650000 508.500000 284.350000 ;
      RECT 416.500000 283.650000 458.500000 284.350000 ;
      RECT 366.500000 283.650000 408.500000 284.350000 ;
      RECT 316.500000 283.650000 358.500000 284.350000 ;
      RECT 266.500000 283.650000 308.500000 284.350000 ;
      RECT 216.500000 283.650000 258.500000 284.350000 ;
      RECT 166.500000 283.650000 208.500000 284.350000 ;
      RECT 116.500000 283.650000 158.500000 284.350000 ;
      RECT 66.500000 283.650000 108.500000 284.350000 ;
      RECT 29.500000 283.650000 58.500000 284.350000 ;
      RECT 0.000000 283.650000 16.500000 284.350000 ;
      RECT 1169.500000 282.350000 1170.500000 283.650000 ;
      RECT 1116.500000 282.350000 1149.500000 283.650000 ;
      RECT 1107.500000 282.350000 1108.500000 283.650000 ;
      RECT 1066.500000 282.350000 1099.500000 283.650000 ;
      RECT 1057.500000 282.350000 1058.500000 283.650000 ;
      RECT 1016.500000 282.350000 1049.500000 283.650000 ;
      RECT 1007.500000 282.350000 1008.500000 283.650000 ;
      RECT 966.500000 282.350000 999.500000 283.650000 ;
      RECT 957.500000 282.350000 958.500000 283.650000 ;
      RECT 916.500000 282.350000 949.500000 283.650000 ;
      RECT 907.500000 282.350000 908.500000 283.650000 ;
      RECT 866.500000 282.350000 899.500000 283.650000 ;
      RECT 857.500000 282.350000 858.500000 283.650000 ;
      RECT 816.500000 282.350000 849.500000 283.650000 ;
      RECT 807.500000 282.350000 808.500000 283.650000 ;
      RECT 766.500000 282.350000 799.500000 283.650000 ;
      RECT 757.500000 282.350000 758.500000 283.650000 ;
      RECT 716.500000 282.350000 749.500000 283.650000 ;
      RECT 707.500000 282.350000 708.500000 283.650000 ;
      RECT 666.500000 282.350000 699.500000 283.650000 ;
      RECT 657.500000 282.350000 658.500000 283.650000 ;
      RECT 616.500000 282.350000 649.500000 283.650000 ;
      RECT 607.500000 282.350000 608.500000 283.650000 ;
      RECT 566.500000 282.350000 599.500000 283.650000 ;
      RECT 557.500000 282.350000 558.500000 283.650000 ;
      RECT 516.500000 282.350000 549.500000 283.650000 ;
      RECT 507.500000 282.350000 508.500000 283.650000 ;
      RECT 466.500000 282.350000 499.500000 283.650000 ;
      RECT 457.500000 282.350000 458.500000 283.650000 ;
      RECT 416.500000 282.350000 449.500000 283.650000 ;
      RECT 407.500000 282.350000 408.500000 283.650000 ;
      RECT 366.500000 282.350000 399.500000 283.650000 ;
      RECT 357.500000 282.350000 358.500000 283.650000 ;
      RECT 316.500000 282.350000 349.500000 283.650000 ;
      RECT 307.500000 282.350000 308.500000 283.650000 ;
      RECT 266.500000 282.350000 299.500000 283.650000 ;
      RECT 257.500000 282.350000 258.500000 283.650000 ;
      RECT 216.500000 282.350000 249.500000 283.650000 ;
      RECT 207.500000 282.350000 208.500000 283.650000 ;
      RECT 166.500000 282.350000 199.500000 283.650000 ;
      RECT 157.500000 282.350000 158.500000 283.650000 ;
      RECT 116.500000 282.350000 149.500000 283.650000 ;
      RECT 107.500000 282.350000 108.500000 283.650000 ;
      RECT 66.500000 282.350000 99.500000 283.650000 ;
      RECT 57.500000 282.350000 58.500000 283.650000 ;
      RECT 29.500000 282.350000 49.500000 283.650000 ;
      RECT 15.500000 282.350000 16.500000 283.650000 ;
      RECT 1157.500000 281.650000 1170.500000 282.350000 ;
      RECT 1107.500000 281.650000 1149.500000 282.350000 ;
      RECT 1057.500000 281.650000 1099.500000 282.350000 ;
      RECT 1007.500000 281.650000 1049.500000 282.350000 ;
      RECT 957.500000 281.650000 999.500000 282.350000 ;
      RECT 907.500000 281.650000 949.500000 282.350000 ;
      RECT 857.500000 281.650000 899.500000 282.350000 ;
      RECT 807.500000 281.650000 849.500000 282.350000 ;
      RECT 757.500000 281.650000 799.500000 282.350000 ;
      RECT 707.500000 281.650000 749.500000 282.350000 ;
      RECT 657.500000 281.650000 699.500000 282.350000 ;
      RECT 607.500000 281.650000 649.500000 282.350000 ;
      RECT 557.500000 281.650000 599.500000 282.350000 ;
      RECT 507.500000 281.650000 549.500000 282.350000 ;
      RECT 457.500000 281.650000 499.500000 282.350000 ;
      RECT 407.500000 281.650000 449.500000 282.350000 ;
      RECT 357.500000 281.650000 399.500000 282.350000 ;
      RECT 307.500000 281.650000 349.500000 282.350000 ;
      RECT 257.500000 281.650000 299.500000 282.350000 ;
      RECT 207.500000 281.650000 249.500000 282.350000 ;
      RECT 157.500000 281.650000 199.500000 282.350000 ;
      RECT 107.500000 281.650000 149.500000 282.350000 ;
      RECT 57.500000 281.650000 99.500000 282.350000 ;
      RECT 15.500000 281.650000 49.500000 282.350000 ;
      RECT 1183.500000 280.350000 1186.000000 283.650000 ;
      RECT 1169.500000 280.350000 1170.500000 281.650000 ;
      RECT 1116.500000 280.350000 1149.500000 281.650000 ;
      RECT 1107.500000 280.350000 1108.500000 281.650000 ;
      RECT 1066.500000 280.350000 1099.500000 281.650000 ;
      RECT 1057.500000 280.350000 1058.500000 281.650000 ;
      RECT 1016.500000 280.350000 1049.500000 281.650000 ;
      RECT 1007.500000 280.350000 1008.500000 281.650000 ;
      RECT 966.500000 280.350000 999.500000 281.650000 ;
      RECT 957.500000 280.350000 958.500000 281.650000 ;
      RECT 916.500000 280.350000 949.500000 281.650000 ;
      RECT 907.500000 280.350000 908.500000 281.650000 ;
      RECT 866.500000 280.350000 899.500000 281.650000 ;
      RECT 857.500000 280.350000 858.500000 281.650000 ;
      RECT 816.500000 280.350000 849.500000 281.650000 ;
      RECT 807.500000 280.350000 808.500000 281.650000 ;
      RECT 766.500000 280.350000 799.500000 281.650000 ;
      RECT 757.500000 280.350000 758.500000 281.650000 ;
      RECT 716.500000 280.350000 749.500000 281.650000 ;
      RECT 707.500000 280.350000 708.500000 281.650000 ;
      RECT 666.500000 280.350000 699.500000 281.650000 ;
      RECT 657.500000 280.350000 658.500000 281.650000 ;
      RECT 616.500000 280.350000 649.500000 281.650000 ;
      RECT 607.500000 280.350000 608.500000 281.650000 ;
      RECT 566.500000 280.350000 599.500000 281.650000 ;
      RECT 557.500000 280.350000 558.500000 281.650000 ;
      RECT 516.500000 280.350000 549.500000 281.650000 ;
      RECT 507.500000 280.350000 508.500000 281.650000 ;
      RECT 466.500000 280.350000 499.500000 281.650000 ;
      RECT 457.500000 280.350000 458.500000 281.650000 ;
      RECT 416.500000 280.350000 449.500000 281.650000 ;
      RECT 407.500000 280.350000 408.500000 281.650000 ;
      RECT 366.500000 280.350000 399.500000 281.650000 ;
      RECT 357.500000 280.350000 358.500000 281.650000 ;
      RECT 316.500000 280.350000 349.500000 281.650000 ;
      RECT 307.500000 280.350000 308.500000 281.650000 ;
      RECT 266.500000 280.350000 299.500000 281.650000 ;
      RECT 257.500000 280.350000 258.500000 281.650000 ;
      RECT 216.500000 280.350000 249.500000 281.650000 ;
      RECT 207.500000 280.350000 208.500000 281.650000 ;
      RECT 166.500000 280.350000 199.500000 281.650000 ;
      RECT 157.500000 280.350000 158.500000 281.650000 ;
      RECT 116.500000 280.350000 149.500000 281.650000 ;
      RECT 107.500000 280.350000 108.500000 281.650000 ;
      RECT 66.500000 280.350000 99.500000 281.650000 ;
      RECT 57.500000 280.350000 58.500000 281.650000 ;
      RECT 29.500000 280.350000 49.500000 281.650000 ;
      RECT 15.500000 280.350000 16.500000 281.650000 ;
      RECT 0.000000 280.350000 2.500000 283.650000 ;
      RECT 1169.500000 279.650000 1186.000000 280.350000 ;
      RECT 1116.500000 279.650000 1156.500000 280.350000 ;
      RECT 1066.500000 279.650000 1108.500000 280.350000 ;
      RECT 1016.500000 279.650000 1058.500000 280.350000 ;
      RECT 966.500000 279.650000 1008.500000 280.350000 ;
      RECT 916.500000 279.650000 958.500000 280.350000 ;
      RECT 866.500000 279.650000 908.500000 280.350000 ;
      RECT 816.500000 279.650000 858.500000 280.350000 ;
      RECT 766.500000 279.650000 808.500000 280.350000 ;
      RECT 716.500000 279.650000 758.500000 280.350000 ;
      RECT 666.500000 279.650000 708.500000 280.350000 ;
      RECT 616.500000 279.650000 658.500000 280.350000 ;
      RECT 566.500000 279.650000 608.500000 280.350000 ;
      RECT 516.500000 279.650000 558.500000 280.350000 ;
      RECT 466.500000 279.650000 508.500000 280.350000 ;
      RECT 416.500000 279.650000 458.500000 280.350000 ;
      RECT 366.500000 279.650000 408.500000 280.350000 ;
      RECT 316.500000 279.650000 358.500000 280.350000 ;
      RECT 266.500000 279.650000 308.500000 280.350000 ;
      RECT 216.500000 279.650000 258.500000 280.350000 ;
      RECT 166.500000 279.650000 208.500000 280.350000 ;
      RECT 116.500000 279.650000 158.500000 280.350000 ;
      RECT 66.500000 279.650000 108.500000 280.350000 ;
      RECT 29.500000 279.650000 58.500000 280.350000 ;
      RECT 0.000000 279.650000 16.500000 280.350000 ;
      RECT 1169.500000 278.350000 1170.500000 279.650000 ;
      RECT 1116.500000 278.350000 1149.500000 279.650000 ;
      RECT 1107.500000 278.350000 1108.500000 279.650000 ;
      RECT 1066.500000 278.350000 1099.500000 279.650000 ;
      RECT 1057.500000 278.350000 1058.500000 279.650000 ;
      RECT 1016.500000 278.350000 1049.500000 279.650000 ;
      RECT 1007.500000 278.350000 1008.500000 279.650000 ;
      RECT 966.500000 278.350000 999.500000 279.650000 ;
      RECT 957.500000 278.350000 958.500000 279.650000 ;
      RECT 916.500000 278.350000 949.500000 279.650000 ;
      RECT 907.500000 278.350000 908.500000 279.650000 ;
      RECT 866.500000 278.350000 899.500000 279.650000 ;
      RECT 857.500000 278.350000 858.500000 279.650000 ;
      RECT 816.500000 278.350000 849.500000 279.650000 ;
      RECT 807.500000 278.350000 808.500000 279.650000 ;
      RECT 766.500000 278.350000 799.500000 279.650000 ;
      RECT 757.500000 278.350000 758.500000 279.650000 ;
      RECT 716.500000 278.350000 749.500000 279.650000 ;
      RECT 707.500000 278.350000 708.500000 279.650000 ;
      RECT 666.500000 278.350000 699.500000 279.650000 ;
      RECT 657.500000 278.350000 658.500000 279.650000 ;
      RECT 616.500000 278.350000 649.500000 279.650000 ;
      RECT 607.500000 278.350000 608.500000 279.650000 ;
      RECT 566.500000 278.350000 599.500000 279.650000 ;
      RECT 557.500000 278.350000 558.500000 279.650000 ;
      RECT 516.500000 278.350000 549.500000 279.650000 ;
      RECT 507.500000 278.350000 508.500000 279.650000 ;
      RECT 466.500000 278.350000 499.500000 279.650000 ;
      RECT 457.500000 278.350000 458.500000 279.650000 ;
      RECT 416.500000 278.350000 449.500000 279.650000 ;
      RECT 407.500000 278.350000 408.500000 279.650000 ;
      RECT 366.500000 278.350000 399.500000 279.650000 ;
      RECT 357.500000 278.350000 358.500000 279.650000 ;
      RECT 316.500000 278.350000 349.500000 279.650000 ;
      RECT 307.500000 278.350000 308.500000 279.650000 ;
      RECT 266.500000 278.350000 299.500000 279.650000 ;
      RECT 257.500000 278.350000 258.500000 279.650000 ;
      RECT 216.500000 278.350000 249.500000 279.650000 ;
      RECT 207.500000 278.350000 208.500000 279.650000 ;
      RECT 166.500000 278.350000 199.500000 279.650000 ;
      RECT 157.500000 278.350000 158.500000 279.650000 ;
      RECT 116.500000 278.350000 149.500000 279.650000 ;
      RECT 107.500000 278.350000 108.500000 279.650000 ;
      RECT 66.500000 278.350000 99.500000 279.650000 ;
      RECT 57.500000 278.350000 58.500000 279.650000 ;
      RECT 29.500000 278.350000 49.500000 279.650000 ;
      RECT 15.500000 278.350000 16.500000 279.650000 ;
      RECT 1157.500000 277.650000 1170.500000 278.350000 ;
      RECT 1107.500000 277.650000 1149.500000 278.350000 ;
      RECT 1057.500000 277.650000 1099.500000 278.350000 ;
      RECT 1007.500000 277.650000 1049.500000 278.350000 ;
      RECT 957.500000 277.650000 999.500000 278.350000 ;
      RECT 907.500000 277.650000 949.500000 278.350000 ;
      RECT 857.500000 277.650000 899.500000 278.350000 ;
      RECT 807.500000 277.650000 849.500000 278.350000 ;
      RECT 757.500000 277.650000 799.500000 278.350000 ;
      RECT 707.500000 277.650000 749.500000 278.350000 ;
      RECT 657.500000 277.650000 699.500000 278.350000 ;
      RECT 607.500000 277.650000 649.500000 278.350000 ;
      RECT 557.500000 277.650000 599.500000 278.350000 ;
      RECT 507.500000 277.650000 549.500000 278.350000 ;
      RECT 457.500000 277.650000 499.500000 278.350000 ;
      RECT 407.500000 277.650000 449.500000 278.350000 ;
      RECT 357.500000 277.650000 399.500000 278.350000 ;
      RECT 307.500000 277.650000 349.500000 278.350000 ;
      RECT 257.500000 277.650000 299.500000 278.350000 ;
      RECT 207.500000 277.650000 249.500000 278.350000 ;
      RECT 157.500000 277.650000 199.500000 278.350000 ;
      RECT 107.500000 277.650000 149.500000 278.350000 ;
      RECT 57.500000 277.650000 99.500000 278.350000 ;
      RECT 15.500000 277.650000 49.500000 278.350000 ;
      RECT 1183.500000 276.350000 1186.000000 279.650000 ;
      RECT 1169.500000 276.350000 1170.500000 277.650000 ;
      RECT 1116.500000 276.350000 1149.500000 277.650000 ;
      RECT 1107.500000 276.350000 1108.500000 277.650000 ;
      RECT 1066.500000 276.350000 1099.500000 277.650000 ;
      RECT 1057.500000 276.350000 1058.500000 277.650000 ;
      RECT 1016.500000 276.350000 1049.500000 277.650000 ;
      RECT 1007.500000 276.350000 1008.500000 277.650000 ;
      RECT 966.500000 276.350000 999.500000 277.650000 ;
      RECT 957.500000 276.350000 958.500000 277.650000 ;
      RECT 916.500000 276.350000 949.500000 277.650000 ;
      RECT 907.500000 276.350000 908.500000 277.650000 ;
      RECT 866.500000 276.350000 899.500000 277.650000 ;
      RECT 857.500000 276.350000 858.500000 277.650000 ;
      RECT 816.500000 276.350000 849.500000 277.650000 ;
      RECT 807.500000 276.350000 808.500000 277.650000 ;
      RECT 766.500000 276.350000 799.500000 277.650000 ;
      RECT 757.500000 276.350000 758.500000 277.650000 ;
      RECT 716.500000 276.350000 749.500000 277.650000 ;
      RECT 707.500000 276.350000 708.500000 277.650000 ;
      RECT 666.500000 276.350000 699.500000 277.650000 ;
      RECT 657.500000 276.350000 658.500000 277.650000 ;
      RECT 616.500000 276.350000 649.500000 277.650000 ;
      RECT 607.500000 276.350000 608.500000 277.650000 ;
      RECT 566.500000 276.350000 599.500000 277.650000 ;
      RECT 557.500000 276.350000 558.500000 277.650000 ;
      RECT 516.500000 276.350000 549.500000 277.650000 ;
      RECT 507.500000 276.350000 508.500000 277.650000 ;
      RECT 466.500000 276.350000 499.500000 277.650000 ;
      RECT 457.500000 276.350000 458.500000 277.650000 ;
      RECT 416.500000 276.350000 449.500000 277.650000 ;
      RECT 407.500000 276.350000 408.500000 277.650000 ;
      RECT 366.500000 276.350000 399.500000 277.650000 ;
      RECT 357.500000 276.350000 358.500000 277.650000 ;
      RECT 316.500000 276.350000 349.500000 277.650000 ;
      RECT 307.500000 276.350000 308.500000 277.650000 ;
      RECT 266.500000 276.350000 299.500000 277.650000 ;
      RECT 257.500000 276.350000 258.500000 277.650000 ;
      RECT 216.500000 276.350000 249.500000 277.650000 ;
      RECT 207.500000 276.350000 208.500000 277.650000 ;
      RECT 166.500000 276.350000 199.500000 277.650000 ;
      RECT 157.500000 276.350000 158.500000 277.650000 ;
      RECT 116.500000 276.350000 149.500000 277.650000 ;
      RECT 107.500000 276.350000 108.500000 277.650000 ;
      RECT 66.500000 276.350000 99.500000 277.650000 ;
      RECT 57.500000 276.350000 58.500000 277.650000 ;
      RECT 29.500000 276.350000 49.500000 277.650000 ;
      RECT 15.500000 276.350000 16.500000 277.650000 ;
      RECT 0.000000 276.350000 2.500000 279.650000 ;
      RECT 1169.500000 275.650000 1186.000000 276.350000 ;
      RECT 1116.500000 275.650000 1156.500000 276.350000 ;
      RECT 1066.500000 275.650000 1108.500000 276.350000 ;
      RECT 1016.500000 275.650000 1058.500000 276.350000 ;
      RECT 966.500000 275.650000 1008.500000 276.350000 ;
      RECT 916.500000 275.650000 958.500000 276.350000 ;
      RECT 866.500000 275.650000 908.500000 276.350000 ;
      RECT 816.500000 275.650000 858.500000 276.350000 ;
      RECT 766.500000 275.650000 808.500000 276.350000 ;
      RECT 716.500000 275.650000 758.500000 276.350000 ;
      RECT 666.500000 275.650000 708.500000 276.350000 ;
      RECT 616.500000 275.650000 658.500000 276.350000 ;
      RECT 566.500000 275.650000 608.500000 276.350000 ;
      RECT 516.500000 275.650000 558.500000 276.350000 ;
      RECT 466.500000 275.650000 508.500000 276.350000 ;
      RECT 416.500000 275.650000 458.500000 276.350000 ;
      RECT 366.500000 275.650000 408.500000 276.350000 ;
      RECT 316.500000 275.650000 358.500000 276.350000 ;
      RECT 266.500000 275.650000 308.500000 276.350000 ;
      RECT 216.500000 275.650000 258.500000 276.350000 ;
      RECT 166.500000 275.650000 208.500000 276.350000 ;
      RECT 116.500000 275.650000 158.500000 276.350000 ;
      RECT 66.500000 275.650000 108.500000 276.350000 ;
      RECT 29.500000 275.650000 58.500000 276.350000 ;
      RECT 0.000000 275.650000 16.500000 276.350000 ;
      RECT 1169.500000 274.350000 1170.500000 275.650000 ;
      RECT 1116.500000 274.350000 1149.500000 275.650000 ;
      RECT 1107.500000 274.350000 1108.500000 275.650000 ;
      RECT 1066.500000 274.350000 1099.500000 275.650000 ;
      RECT 1057.500000 274.350000 1058.500000 275.650000 ;
      RECT 1016.500000 274.350000 1049.500000 275.650000 ;
      RECT 1007.500000 274.350000 1008.500000 275.650000 ;
      RECT 966.500000 274.350000 999.500000 275.650000 ;
      RECT 957.500000 274.350000 958.500000 275.650000 ;
      RECT 916.500000 274.350000 949.500000 275.650000 ;
      RECT 907.500000 274.350000 908.500000 275.650000 ;
      RECT 866.500000 274.350000 899.500000 275.650000 ;
      RECT 857.500000 274.350000 858.500000 275.650000 ;
      RECT 816.500000 274.350000 849.500000 275.650000 ;
      RECT 807.500000 274.350000 808.500000 275.650000 ;
      RECT 766.500000 274.350000 799.500000 275.650000 ;
      RECT 757.500000 274.350000 758.500000 275.650000 ;
      RECT 716.500000 274.350000 749.500000 275.650000 ;
      RECT 707.500000 274.350000 708.500000 275.650000 ;
      RECT 666.500000 274.350000 699.500000 275.650000 ;
      RECT 657.500000 274.350000 658.500000 275.650000 ;
      RECT 616.500000 274.350000 649.500000 275.650000 ;
      RECT 607.500000 274.350000 608.500000 275.650000 ;
      RECT 566.500000 274.350000 599.500000 275.650000 ;
      RECT 557.500000 274.350000 558.500000 275.650000 ;
      RECT 516.500000 274.350000 549.500000 275.650000 ;
      RECT 507.500000 274.350000 508.500000 275.650000 ;
      RECT 466.500000 274.350000 499.500000 275.650000 ;
      RECT 457.500000 274.350000 458.500000 275.650000 ;
      RECT 416.500000 274.350000 449.500000 275.650000 ;
      RECT 407.500000 274.350000 408.500000 275.650000 ;
      RECT 366.500000 274.350000 399.500000 275.650000 ;
      RECT 357.500000 274.350000 358.500000 275.650000 ;
      RECT 316.500000 274.350000 349.500000 275.650000 ;
      RECT 307.500000 274.350000 308.500000 275.650000 ;
      RECT 266.500000 274.350000 299.500000 275.650000 ;
      RECT 257.500000 274.350000 258.500000 275.650000 ;
      RECT 216.500000 274.350000 249.500000 275.650000 ;
      RECT 207.500000 274.350000 208.500000 275.650000 ;
      RECT 166.500000 274.350000 199.500000 275.650000 ;
      RECT 157.500000 274.350000 158.500000 275.650000 ;
      RECT 116.500000 274.350000 149.500000 275.650000 ;
      RECT 107.500000 274.350000 108.500000 275.650000 ;
      RECT 66.500000 274.350000 99.500000 275.650000 ;
      RECT 57.500000 274.350000 58.500000 275.650000 ;
      RECT 29.500000 274.350000 49.500000 275.650000 ;
      RECT 15.500000 274.350000 16.500000 275.650000 ;
      RECT 1157.500000 273.650000 1170.500000 274.350000 ;
      RECT 1107.500000 273.650000 1149.500000 274.350000 ;
      RECT 1057.500000 273.650000 1099.500000 274.350000 ;
      RECT 1007.500000 273.650000 1049.500000 274.350000 ;
      RECT 957.500000 273.650000 999.500000 274.350000 ;
      RECT 907.500000 273.650000 949.500000 274.350000 ;
      RECT 857.500000 273.650000 899.500000 274.350000 ;
      RECT 807.500000 273.650000 849.500000 274.350000 ;
      RECT 757.500000 273.650000 799.500000 274.350000 ;
      RECT 707.500000 273.650000 749.500000 274.350000 ;
      RECT 657.500000 273.650000 699.500000 274.350000 ;
      RECT 607.500000 273.650000 649.500000 274.350000 ;
      RECT 557.500000 273.650000 599.500000 274.350000 ;
      RECT 507.500000 273.650000 549.500000 274.350000 ;
      RECT 457.500000 273.650000 499.500000 274.350000 ;
      RECT 407.500000 273.650000 449.500000 274.350000 ;
      RECT 357.500000 273.650000 399.500000 274.350000 ;
      RECT 307.500000 273.650000 349.500000 274.350000 ;
      RECT 257.500000 273.650000 299.500000 274.350000 ;
      RECT 207.500000 273.650000 249.500000 274.350000 ;
      RECT 157.500000 273.650000 199.500000 274.350000 ;
      RECT 107.500000 273.650000 149.500000 274.350000 ;
      RECT 57.500000 273.650000 99.500000 274.350000 ;
      RECT 15.500000 273.650000 49.500000 274.350000 ;
      RECT 1183.500000 272.350000 1186.000000 275.650000 ;
      RECT 1169.500000 272.350000 1170.500000 273.650000 ;
      RECT 1116.500000 272.350000 1149.500000 273.650000 ;
      RECT 1107.500000 272.350000 1108.500000 273.650000 ;
      RECT 1066.500000 272.350000 1099.500000 273.650000 ;
      RECT 1057.500000 272.350000 1058.500000 273.650000 ;
      RECT 1016.500000 272.350000 1049.500000 273.650000 ;
      RECT 1007.500000 272.350000 1008.500000 273.650000 ;
      RECT 966.500000 272.350000 999.500000 273.650000 ;
      RECT 957.500000 272.350000 958.500000 273.650000 ;
      RECT 916.500000 272.350000 949.500000 273.650000 ;
      RECT 907.500000 272.350000 908.500000 273.650000 ;
      RECT 866.500000 272.350000 899.500000 273.650000 ;
      RECT 857.500000 272.350000 858.500000 273.650000 ;
      RECT 816.500000 272.350000 849.500000 273.650000 ;
      RECT 807.500000 272.350000 808.500000 273.650000 ;
      RECT 766.500000 272.350000 799.500000 273.650000 ;
      RECT 757.500000 272.350000 758.500000 273.650000 ;
      RECT 716.500000 272.350000 749.500000 273.650000 ;
      RECT 707.500000 272.350000 708.500000 273.650000 ;
      RECT 666.500000 272.350000 699.500000 273.650000 ;
      RECT 657.500000 272.350000 658.500000 273.650000 ;
      RECT 616.500000 272.350000 649.500000 273.650000 ;
      RECT 607.500000 272.350000 608.500000 273.650000 ;
      RECT 566.500000 272.350000 599.500000 273.650000 ;
      RECT 557.500000 272.350000 558.500000 273.650000 ;
      RECT 516.500000 272.350000 549.500000 273.650000 ;
      RECT 507.500000 272.350000 508.500000 273.650000 ;
      RECT 466.500000 272.350000 499.500000 273.650000 ;
      RECT 457.500000 272.350000 458.500000 273.650000 ;
      RECT 416.500000 272.350000 449.500000 273.650000 ;
      RECT 407.500000 272.350000 408.500000 273.650000 ;
      RECT 366.500000 272.350000 399.500000 273.650000 ;
      RECT 357.500000 272.350000 358.500000 273.650000 ;
      RECT 316.500000 272.350000 349.500000 273.650000 ;
      RECT 307.500000 272.350000 308.500000 273.650000 ;
      RECT 266.500000 272.350000 299.500000 273.650000 ;
      RECT 257.500000 272.350000 258.500000 273.650000 ;
      RECT 216.500000 272.350000 249.500000 273.650000 ;
      RECT 207.500000 272.350000 208.500000 273.650000 ;
      RECT 166.500000 272.350000 199.500000 273.650000 ;
      RECT 157.500000 272.350000 158.500000 273.650000 ;
      RECT 116.500000 272.350000 149.500000 273.650000 ;
      RECT 107.500000 272.350000 108.500000 273.650000 ;
      RECT 66.500000 272.350000 99.500000 273.650000 ;
      RECT 57.500000 272.350000 58.500000 273.650000 ;
      RECT 29.500000 272.350000 49.500000 273.650000 ;
      RECT 15.500000 272.350000 16.500000 273.650000 ;
      RECT 0.000000 272.350000 2.500000 275.650000 ;
      RECT 1169.500000 271.650000 1186.000000 272.350000 ;
      RECT 1116.500000 271.650000 1156.500000 272.350000 ;
      RECT 1066.500000 271.650000 1108.500000 272.350000 ;
      RECT 1016.500000 271.650000 1058.500000 272.350000 ;
      RECT 966.500000 271.650000 1008.500000 272.350000 ;
      RECT 916.500000 271.650000 958.500000 272.350000 ;
      RECT 866.500000 271.650000 908.500000 272.350000 ;
      RECT 816.500000 271.650000 858.500000 272.350000 ;
      RECT 766.500000 271.650000 808.500000 272.350000 ;
      RECT 716.500000 271.650000 758.500000 272.350000 ;
      RECT 666.500000 271.650000 708.500000 272.350000 ;
      RECT 616.500000 271.650000 658.500000 272.350000 ;
      RECT 566.500000 271.650000 608.500000 272.350000 ;
      RECT 516.500000 271.650000 558.500000 272.350000 ;
      RECT 466.500000 271.650000 508.500000 272.350000 ;
      RECT 416.500000 271.650000 458.500000 272.350000 ;
      RECT 366.500000 271.650000 408.500000 272.350000 ;
      RECT 316.500000 271.650000 358.500000 272.350000 ;
      RECT 266.500000 271.650000 308.500000 272.350000 ;
      RECT 216.500000 271.650000 258.500000 272.350000 ;
      RECT 166.500000 271.650000 208.500000 272.350000 ;
      RECT 116.500000 271.650000 158.500000 272.350000 ;
      RECT 66.500000 271.650000 108.500000 272.350000 ;
      RECT 29.500000 271.650000 58.500000 272.350000 ;
      RECT 0.000000 271.650000 16.500000 272.350000 ;
      RECT 1169.500000 270.350000 1170.500000 271.650000 ;
      RECT 1116.500000 270.350000 1149.500000 271.650000 ;
      RECT 1107.500000 270.350000 1108.500000 271.650000 ;
      RECT 1066.500000 270.350000 1099.500000 271.650000 ;
      RECT 1057.500000 270.350000 1058.500000 271.650000 ;
      RECT 1016.500000 270.350000 1049.500000 271.650000 ;
      RECT 1007.500000 270.350000 1008.500000 271.650000 ;
      RECT 966.500000 270.350000 999.500000 271.650000 ;
      RECT 957.500000 270.350000 958.500000 271.650000 ;
      RECT 916.500000 270.350000 949.500000 271.650000 ;
      RECT 907.500000 270.350000 908.500000 271.650000 ;
      RECT 866.500000 270.350000 899.500000 271.650000 ;
      RECT 857.500000 270.350000 858.500000 271.650000 ;
      RECT 816.500000 270.350000 849.500000 271.650000 ;
      RECT 807.500000 270.350000 808.500000 271.650000 ;
      RECT 766.500000 270.350000 799.500000 271.650000 ;
      RECT 757.500000 270.350000 758.500000 271.650000 ;
      RECT 716.500000 270.350000 749.500000 271.650000 ;
      RECT 707.500000 270.350000 708.500000 271.650000 ;
      RECT 666.500000 270.350000 699.500000 271.650000 ;
      RECT 657.500000 270.350000 658.500000 271.650000 ;
      RECT 616.500000 270.350000 649.500000 271.650000 ;
      RECT 607.500000 270.350000 608.500000 271.650000 ;
      RECT 566.500000 270.350000 599.500000 271.650000 ;
      RECT 557.500000 270.350000 558.500000 271.650000 ;
      RECT 516.500000 270.350000 549.500000 271.650000 ;
      RECT 507.500000 270.350000 508.500000 271.650000 ;
      RECT 466.500000 270.350000 499.500000 271.650000 ;
      RECT 457.500000 270.350000 458.500000 271.650000 ;
      RECT 416.500000 270.350000 449.500000 271.650000 ;
      RECT 407.500000 270.350000 408.500000 271.650000 ;
      RECT 366.500000 270.350000 399.500000 271.650000 ;
      RECT 357.500000 270.350000 358.500000 271.650000 ;
      RECT 316.500000 270.350000 349.500000 271.650000 ;
      RECT 307.500000 270.350000 308.500000 271.650000 ;
      RECT 266.500000 270.350000 299.500000 271.650000 ;
      RECT 257.500000 270.350000 258.500000 271.650000 ;
      RECT 216.500000 270.350000 249.500000 271.650000 ;
      RECT 207.500000 270.350000 208.500000 271.650000 ;
      RECT 166.500000 270.350000 199.500000 271.650000 ;
      RECT 157.500000 270.350000 158.500000 271.650000 ;
      RECT 116.500000 270.350000 149.500000 271.650000 ;
      RECT 107.500000 270.350000 108.500000 271.650000 ;
      RECT 66.500000 270.350000 99.500000 271.650000 ;
      RECT 57.500000 270.350000 58.500000 271.650000 ;
      RECT 29.500000 270.350000 49.500000 271.650000 ;
      RECT 15.500000 270.350000 16.500000 271.650000 ;
      RECT 1157.500000 269.650000 1170.500000 270.350000 ;
      RECT 1107.500000 269.650000 1149.500000 270.350000 ;
      RECT 1057.500000 269.650000 1099.500000 270.350000 ;
      RECT 1007.500000 269.650000 1049.500000 270.350000 ;
      RECT 957.500000 269.650000 999.500000 270.350000 ;
      RECT 907.500000 269.650000 949.500000 270.350000 ;
      RECT 857.500000 269.650000 899.500000 270.350000 ;
      RECT 807.500000 269.650000 849.500000 270.350000 ;
      RECT 757.500000 269.650000 799.500000 270.350000 ;
      RECT 707.500000 269.650000 749.500000 270.350000 ;
      RECT 657.500000 269.650000 699.500000 270.350000 ;
      RECT 607.500000 269.650000 649.500000 270.350000 ;
      RECT 557.500000 269.650000 599.500000 270.350000 ;
      RECT 507.500000 269.650000 549.500000 270.350000 ;
      RECT 457.500000 269.650000 499.500000 270.350000 ;
      RECT 407.500000 269.650000 449.500000 270.350000 ;
      RECT 357.500000 269.650000 399.500000 270.350000 ;
      RECT 307.500000 269.650000 349.500000 270.350000 ;
      RECT 257.500000 269.650000 299.500000 270.350000 ;
      RECT 207.500000 269.650000 249.500000 270.350000 ;
      RECT 157.500000 269.650000 199.500000 270.350000 ;
      RECT 107.500000 269.650000 149.500000 270.350000 ;
      RECT 57.500000 269.650000 99.500000 270.350000 ;
      RECT 15.500000 269.650000 49.500000 270.350000 ;
      RECT 1183.500000 268.350000 1186.000000 271.650000 ;
      RECT 1169.500000 268.350000 1170.500000 269.650000 ;
      RECT 1116.500000 268.350000 1149.500000 269.650000 ;
      RECT 1107.500000 268.350000 1108.500000 269.650000 ;
      RECT 1066.500000 268.350000 1099.500000 269.650000 ;
      RECT 1057.500000 268.350000 1058.500000 269.650000 ;
      RECT 1016.500000 268.350000 1049.500000 269.650000 ;
      RECT 1007.500000 268.350000 1008.500000 269.650000 ;
      RECT 966.500000 268.350000 999.500000 269.650000 ;
      RECT 957.500000 268.350000 958.500000 269.650000 ;
      RECT 916.500000 268.350000 949.500000 269.650000 ;
      RECT 907.500000 268.350000 908.500000 269.650000 ;
      RECT 866.500000 268.350000 899.500000 269.650000 ;
      RECT 857.500000 268.350000 858.500000 269.650000 ;
      RECT 816.500000 268.350000 849.500000 269.650000 ;
      RECT 807.500000 268.350000 808.500000 269.650000 ;
      RECT 766.500000 268.350000 799.500000 269.650000 ;
      RECT 757.500000 268.350000 758.500000 269.650000 ;
      RECT 716.500000 268.350000 749.500000 269.650000 ;
      RECT 707.500000 268.350000 708.500000 269.650000 ;
      RECT 666.500000 268.350000 699.500000 269.650000 ;
      RECT 657.500000 268.350000 658.500000 269.650000 ;
      RECT 616.500000 268.350000 649.500000 269.650000 ;
      RECT 607.500000 268.350000 608.500000 269.650000 ;
      RECT 566.500000 268.350000 599.500000 269.650000 ;
      RECT 557.500000 268.350000 558.500000 269.650000 ;
      RECT 516.500000 268.350000 549.500000 269.650000 ;
      RECT 507.500000 268.350000 508.500000 269.650000 ;
      RECT 466.500000 268.350000 499.500000 269.650000 ;
      RECT 457.500000 268.350000 458.500000 269.650000 ;
      RECT 416.500000 268.350000 449.500000 269.650000 ;
      RECT 407.500000 268.350000 408.500000 269.650000 ;
      RECT 366.500000 268.350000 399.500000 269.650000 ;
      RECT 357.500000 268.350000 358.500000 269.650000 ;
      RECT 316.500000 268.350000 349.500000 269.650000 ;
      RECT 307.500000 268.350000 308.500000 269.650000 ;
      RECT 266.500000 268.350000 299.500000 269.650000 ;
      RECT 257.500000 268.350000 258.500000 269.650000 ;
      RECT 216.500000 268.350000 249.500000 269.650000 ;
      RECT 207.500000 268.350000 208.500000 269.650000 ;
      RECT 166.500000 268.350000 199.500000 269.650000 ;
      RECT 157.500000 268.350000 158.500000 269.650000 ;
      RECT 116.500000 268.350000 149.500000 269.650000 ;
      RECT 107.500000 268.350000 108.500000 269.650000 ;
      RECT 66.500000 268.350000 99.500000 269.650000 ;
      RECT 57.500000 268.350000 58.500000 269.650000 ;
      RECT 29.500000 268.350000 49.500000 269.650000 ;
      RECT 15.500000 268.350000 16.500000 269.650000 ;
      RECT 0.000000 268.350000 2.500000 271.650000 ;
      RECT 1169.500000 267.650000 1186.000000 268.350000 ;
      RECT 1116.500000 267.650000 1156.500000 268.350000 ;
      RECT 1066.500000 267.650000 1108.500000 268.350000 ;
      RECT 1016.500000 267.650000 1058.500000 268.350000 ;
      RECT 966.500000 267.650000 1008.500000 268.350000 ;
      RECT 916.500000 267.650000 958.500000 268.350000 ;
      RECT 866.500000 267.650000 908.500000 268.350000 ;
      RECT 816.500000 267.650000 858.500000 268.350000 ;
      RECT 766.500000 267.650000 808.500000 268.350000 ;
      RECT 716.500000 267.650000 758.500000 268.350000 ;
      RECT 666.500000 267.650000 708.500000 268.350000 ;
      RECT 616.500000 267.650000 658.500000 268.350000 ;
      RECT 566.500000 267.650000 608.500000 268.350000 ;
      RECT 516.500000 267.650000 558.500000 268.350000 ;
      RECT 466.500000 267.650000 508.500000 268.350000 ;
      RECT 416.500000 267.650000 458.500000 268.350000 ;
      RECT 366.500000 267.650000 408.500000 268.350000 ;
      RECT 316.500000 267.650000 358.500000 268.350000 ;
      RECT 266.500000 267.650000 308.500000 268.350000 ;
      RECT 216.500000 267.650000 258.500000 268.350000 ;
      RECT 166.500000 267.650000 208.500000 268.350000 ;
      RECT 116.500000 267.650000 158.500000 268.350000 ;
      RECT 66.500000 267.650000 108.500000 268.350000 ;
      RECT 29.500000 267.650000 58.500000 268.350000 ;
      RECT 0.000000 267.650000 16.500000 268.350000 ;
      RECT 1169.500000 266.350000 1170.500000 267.650000 ;
      RECT 1116.500000 266.350000 1149.500000 267.650000 ;
      RECT 1107.500000 266.350000 1108.500000 267.650000 ;
      RECT 1066.500000 266.350000 1099.500000 267.650000 ;
      RECT 1057.500000 266.350000 1058.500000 267.650000 ;
      RECT 1016.500000 266.350000 1049.500000 267.650000 ;
      RECT 1007.500000 266.350000 1008.500000 267.650000 ;
      RECT 966.500000 266.350000 999.500000 267.650000 ;
      RECT 957.500000 266.350000 958.500000 267.650000 ;
      RECT 916.500000 266.350000 949.500000 267.650000 ;
      RECT 907.500000 266.350000 908.500000 267.650000 ;
      RECT 866.500000 266.350000 899.500000 267.650000 ;
      RECT 857.500000 266.350000 858.500000 267.650000 ;
      RECT 816.500000 266.350000 849.500000 267.650000 ;
      RECT 807.500000 266.350000 808.500000 267.650000 ;
      RECT 766.500000 266.350000 799.500000 267.650000 ;
      RECT 757.500000 266.350000 758.500000 267.650000 ;
      RECT 716.500000 266.350000 749.500000 267.650000 ;
      RECT 707.500000 266.350000 708.500000 267.650000 ;
      RECT 666.500000 266.350000 699.500000 267.650000 ;
      RECT 657.500000 266.350000 658.500000 267.650000 ;
      RECT 616.500000 266.350000 649.500000 267.650000 ;
      RECT 607.500000 266.350000 608.500000 267.650000 ;
      RECT 566.500000 266.350000 599.500000 267.650000 ;
      RECT 557.500000 266.350000 558.500000 267.650000 ;
      RECT 516.500000 266.350000 549.500000 267.650000 ;
      RECT 507.500000 266.350000 508.500000 267.650000 ;
      RECT 466.500000 266.350000 499.500000 267.650000 ;
      RECT 457.500000 266.350000 458.500000 267.650000 ;
      RECT 416.500000 266.350000 449.500000 267.650000 ;
      RECT 407.500000 266.350000 408.500000 267.650000 ;
      RECT 366.500000 266.350000 399.500000 267.650000 ;
      RECT 357.500000 266.350000 358.500000 267.650000 ;
      RECT 316.500000 266.350000 349.500000 267.650000 ;
      RECT 307.500000 266.350000 308.500000 267.650000 ;
      RECT 266.500000 266.350000 299.500000 267.650000 ;
      RECT 257.500000 266.350000 258.500000 267.650000 ;
      RECT 216.500000 266.350000 249.500000 267.650000 ;
      RECT 207.500000 266.350000 208.500000 267.650000 ;
      RECT 166.500000 266.350000 199.500000 267.650000 ;
      RECT 157.500000 266.350000 158.500000 267.650000 ;
      RECT 116.500000 266.350000 149.500000 267.650000 ;
      RECT 107.500000 266.350000 108.500000 267.650000 ;
      RECT 66.500000 266.350000 99.500000 267.650000 ;
      RECT 57.500000 266.350000 58.500000 267.650000 ;
      RECT 29.500000 266.350000 49.500000 267.650000 ;
      RECT 15.500000 266.350000 16.500000 267.650000 ;
      RECT 1157.500000 265.650000 1170.500000 266.350000 ;
      RECT 1107.500000 265.650000 1149.500000 266.350000 ;
      RECT 1057.500000 265.650000 1099.500000 266.350000 ;
      RECT 1007.500000 265.650000 1049.500000 266.350000 ;
      RECT 957.500000 265.650000 999.500000 266.350000 ;
      RECT 907.500000 265.650000 949.500000 266.350000 ;
      RECT 857.500000 265.650000 899.500000 266.350000 ;
      RECT 807.500000 265.650000 849.500000 266.350000 ;
      RECT 757.500000 265.650000 799.500000 266.350000 ;
      RECT 707.500000 265.650000 749.500000 266.350000 ;
      RECT 657.500000 265.650000 699.500000 266.350000 ;
      RECT 607.500000 265.650000 649.500000 266.350000 ;
      RECT 557.500000 265.650000 599.500000 266.350000 ;
      RECT 507.500000 265.650000 549.500000 266.350000 ;
      RECT 457.500000 265.650000 499.500000 266.350000 ;
      RECT 407.500000 265.650000 449.500000 266.350000 ;
      RECT 357.500000 265.650000 399.500000 266.350000 ;
      RECT 307.500000 265.650000 349.500000 266.350000 ;
      RECT 257.500000 265.650000 299.500000 266.350000 ;
      RECT 207.500000 265.650000 249.500000 266.350000 ;
      RECT 157.500000 265.650000 199.500000 266.350000 ;
      RECT 107.500000 265.650000 149.500000 266.350000 ;
      RECT 57.500000 265.650000 99.500000 266.350000 ;
      RECT 15.500000 265.650000 49.500000 266.350000 ;
      RECT 1183.500000 264.350000 1186.000000 267.650000 ;
      RECT 1169.500000 264.350000 1170.500000 265.650000 ;
      RECT 1116.500000 264.350000 1149.500000 265.650000 ;
      RECT 1107.500000 264.350000 1108.500000 265.650000 ;
      RECT 1066.500000 264.350000 1099.500000 265.650000 ;
      RECT 1057.500000 264.350000 1058.500000 265.650000 ;
      RECT 1016.500000 264.350000 1049.500000 265.650000 ;
      RECT 1007.500000 264.350000 1008.500000 265.650000 ;
      RECT 966.500000 264.350000 999.500000 265.650000 ;
      RECT 957.500000 264.350000 958.500000 265.650000 ;
      RECT 916.500000 264.350000 949.500000 265.650000 ;
      RECT 907.500000 264.350000 908.500000 265.650000 ;
      RECT 866.500000 264.350000 899.500000 265.650000 ;
      RECT 857.500000 264.350000 858.500000 265.650000 ;
      RECT 816.500000 264.350000 849.500000 265.650000 ;
      RECT 807.500000 264.350000 808.500000 265.650000 ;
      RECT 766.500000 264.350000 799.500000 265.650000 ;
      RECT 757.500000 264.350000 758.500000 265.650000 ;
      RECT 716.500000 264.350000 749.500000 265.650000 ;
      RECT 707.500000 264.350000 708.500000 265.650000 ;
      RECT 666.500000 264.350000 699.500000 265.650000 ;
      RECT 657.500000 264.350000 658.500000 265.650000 ;
      RECT 616.500000 264.350000 649.500000 265.650000 ;
      RECT 607.500000 264.350000 608.500000 265.650000 ;
      RECT 566.500000 264.350000 599.500000 265.650000 ;
      RECT 557.500000 264.350000 558.500000 265.650000 ;
      RECT 516.500000 264.350000 549.500000 265.650000 ;
      RECT 507.500000 264.350000 508.500000 265.650000 ;
      RECT 466.500000 264.350000 499.500000 265.650000 ;
      RECT 457.500000 264.350000 458.500000 265.650000 ;
      RECT 416.500000 264.350000 449.500000 265.650000 ;
      RECT 407.500000 264.350000 408.500000 265.650000 ;
      RECT 366.500000 264.350000 399.500000 265.650000 ;
      RECT 357.500000 264.350000 358.500000 265.650000 ;
      RECT 316.500000 264.350000 349.500000 265.650000 ;
      RECT 307.500000 264.350000 308.500000 265.650000 ;
      RECT 266.500000 264.350000 299.500000 265.650000 ;
      RECT 257.500000 264.350000 258.500000 265.650000 ;
      RECT 216.500000 264.350000 249.500000 265.650000 ;
      RECT 207.500000 264.350000 208.500000 265.650000 ;
      RECT 166.500000 264.350000 199.500000 265.650000 ;
      RECT 157.500000 264.350000 158.500000 265.650000 ;
      RECT 116.500000 264.350000 149.500000 265.650000 ;
      RECT 107.500000 264.350000 108.500000 265.650000 ;
      RECT 66.500000 264.350000 99.500000 265.650000 ;
      RECT 57.500000 264.350000 58.500000 265.650000 ;
      RECT 29.500000 264.350000 49.500000 265.650000 ;
      RECT 15.500000 264.350000 16.500000 265.650000 ;
      RECT 0.000000 264.350000 2.500000 267.650000 ;
      RECT 1169.500000 263.650000 1186.000000 264.350000 ;
      RECT 1116.500000 263.650000 1156.500000 264.350000 ;
      RECT 1066.500000 263.650000 1108.500000 264.350000 ;
      RECT 1016.500000 263.650000 1058.500000 264.350000 ;
      RECT 966.500000 263.650000 1008.500000 264.350000 ;
      RECT 916.500000 263.650000 958.500000 264.350000 ;
      RECT 866.500000 263.650000 908.500000 264.350000 ;
      RECT 816.500000 263.650000 858.500000 264.350000 ;
      RECT 766.500000 263.650000 808.500000 264.350000 ;
      RECT 716.500000 263.650000 758.500000 264.350000 ;
      RECT 666.500000 263.650000 708.500000 264.350000 ;
      RECT 616.500000 263.650000 658.500000 264.350000 ;
      RECT 566.500000 263.650000 608.500000 264.350000 ;
      RECT 516.500000 263.650000 558.500000 264.350000 ;
      RECT 466.500000 263.650000 508.500000 264.350000 ;
      RECT 416.500000 263.650000 458.500000 264.350000 ;
      RECT 366.500000 263.650000 408.500000 264.350000 ;
      RECT 316.500000 263.650000 358.500000 264.350000 ;
      RECT 266.500000 263.650000 308.500000 264.350000 ;
      RECT 216.500000 263.650000 258.500000 264.350000 ;
      RECT 166.500000 263.650000 208.500000 264.350000 ;
      RECT 116.500000 263.650000 158.500000 264.350000 ;
      RECT 66.500000 263.650000 108.500000 264.350000 ;
      RECT 29.500000 263.650000 58.500000 264.350000 ;
      RECT 0.000000 263.650000 16.500000 264.350000 ;
      RECT 1169.500000 262.350000 1170.500000 263.650000 ;
      RECT 1116.500000 262.350000 1149.500000 263.650000 ;
      RECT 1107.500000 262.350000 1108.500000 263.650000 ;
      RECT 1066.500000 262.350000 1099.500000 263.650000 ;
      RECT 1057.500000 262.350000 1058.500000 263.650000 ;
      RECT 1016.500000 262.350000 1049.500000 263.650000 ;
      RECT 1007.500000 262.350000 1008.500000 263.650000 ;
      RECT 966.500000 262.350000 999.500000 263.650000 ;
      RECT 957.500000 262.350000 958.500000 263.650000 ;
      RECT 916.500000 262.350000 949.500000 263.650000 ;
      RECT 907.500000 262.350000 908.500000 263.650000 ;
      RECT 866.500000 262.350000 899.500000 263.650000 ;
      RECT 857.500000 262.350000 858.500000 263.650000 ;
      RECT 816.500000 262.350000 849.500000 263.650000 ;
      RECT 807.500000 262.350000 808.500000 263.650000 ;
      RECT 766.500000 262.350000 799.500000 263.650000 ;
      RECT 757.500000 262.350000 758.500000 263.650000 ;
      RECT 716.500000 262.350000 749.500000 263.650000 ;
      RECT 707.500000 262.350000 708.500000 263.650000 ;
      RECT 666.500000 262.350000 699.500000 263.650000 ;
      RECT 657.500000 262.350000 658.500000 263.650000 ;
      RECT 616.500000 262.350000 649.500000 263.650000 ;
      RECT 607.500000 262.350000 608.500000 263.650000 ;
      RECT 566.500000 262.350000 599.500000 263.650000 ;
      RECT 557.500000 262.350000 558.500000 263.650000 ;
      RECT 516.500000 262.350000 549.500000 263.650000 ;
      RECT 507.500000 262.350000 508.500000 263.650000 ;
      RECT 466.500000 262.350000 499.500000 263.650000 ;
      RECT 457.500000 262.350000 458.500000 263.650000 ;
      RECT 416.500000 262.350000 449.500000 263.650000 ;
      RECT 407.500000 262.350000 408.500000 263.650000 ;
      RECT 366.500000 262.350000 399.500000 263.650000 ;
      RECT 357.500000 262.350000 358.500000 263.650000 ;
      RECT 316.500000 262.350000 349.500000 263.650000 ;
      RECT 307.500000 262.350000 308.500000 263.650000 ;
      RECT 266.500000 262.350000 299.500000 263.650000 ;
      RECT 257.500000 262.350000 258.500000 263.650000 ;
      RECT 216.500000 262.350000 249.500000 263.650000 ;
      RECT 207.500000 262.350000 208.500000 263.650000 ;
      RECT 166.500000 262.350000 199.500000 263.650000 ;
      RECT 157.500000 262.350000 158.500000 263.650000 ;
      RECT 116.500000 262.350000 149.500000 263.650000 ;
      RECT 107.500000 262.350000 108.500000 263.650000 ;
      RECT 66.500000 262.350000 99.500000 263.650000 ;
      RECT 57.500000 262.350000 58.500000 263.650000 ;
      RECT 29.500000 262.350000 49.500000 263.650000 ;
      RECT 15.500000 262.350000 16.500000 263.650000 ;
      RECT 1157.500000 261.650000 1170.500000 262.350000 ;
      RECT 1107.500000 261.650000 1149.500000 262.350000 ;
      RECT 1057.500000 261.650000 1099.500000 262.350000 ;
      RECT 1007.500000 261.650000 1049.500000 262.350000 ;
      RECT 957.500000 261.650000 999.500000 262.350000 ;
      RECT 907.500000 261.650000 949.500000 262.350000 ;
      RECT 857.500000 261.650000 899.500000 262.350000 ;
      RECT 807.500000 261.650000 849.500000 262.350000 ;
      RECT 757.500000 261.650000 799.500000 262.350000 ;
      RECT 707.500000 261.650000 749.500000 262.350000 ;
      RECT 657.500000 261.650000 699.500000 262.350000 ;
      RECT 607.500000 261.650000 649.500000 262.350000 ;
      RECT 557.500000 261.650000 599.500000 262.350000 ;
      RECT 507.500000 261.650000 549.500000 262.350000 ;
      RECT 457.500000 261.650000 499.500000 262.350000 ;
      RECT 407.500000 261.650000 449.500000 262.350000 ;
      RECT 357.500000 261.650000 399.500000 262.350000 ;
      RECT 307.500000 261.650000 349.500000 262.350000 ;
      RECT 257.500000 261.650000 299.500000 262.350000 ;
      RECT 207.500000 261.650000 249.500000 262.350000 ;
      RECT 157.500000 261.650000 199.500000 262.350000 ;
      RECT 107.500000 261.650000 149.500000 262.350000 ;
      RECT 57.500000 261.650000 99.500000 262.350000 ;
      RECT 15.500000 261.650000 49.500000 262.350000 ;
      RECT 1183.500000 260.350000 1186.000000 263.650000 ;
      RECT 1169.500000 260.350000 1170.500000 261.650000 ;
      RECT 1116.500000 260.350000 1149.500000 261.650000 ;
      RECT 1107.500000 260.350000 1108.500000 261.650000 ;
      RECT 1066.500000 260.350000 1099.500000 261.650000 ;
      RECT 1057.500000 260.350000 1058.500000 261.650000 ;
      RECT 1016.500000 260.350000 1049.500000 261.650000 ;
      RECT 1007.500000 260.350000 1008.500000 261.650000 ;
      RECT 966.500000 260.350000 999.500000 261.650000 ;
      RECT 957.500000 260.350000 958.500000 261.650000 ;
      RECT 916.500000 260.350000 949.500000 261.650000 ;
      RECT 907.500000 260.350000 908.500000 261.650000 ;
      RECT 866.500000 260.350000 899.500000 261.650000 ;
      RECT 857.500000 260.350000 858.500000 261.650000 ;
      RECT 816.500000 260.350000 849.500000 261.650000 ;
      RECT 807.500000 260.350000 808.500000 261.650000 ;
      RECT 766.500000 260.350000 799.500000 261.650000 ;
      RECT 757.500000 260.350000 758.500000 261.650000 ;
      RECT 716.500000 260.350000 749.500000 261.650000 ;
      RECT 707.500000 260.350000 708.500000 261.650000 ;
      RECT 666.500000 260.350000 699.500000 261.650000 ;
      RECT 657.500000 260.350000 658.500000 261.650000 ;
      RECT 616.500000 260.350000 649.500000 261.650000 ;
      RECT 607.500000 260.350000 608.500000 261.650000 ;
      RECT 566.500000 260.350000 599.500000 261.650000 ;
      RECT 557.500000 260.350000 558.500000 261.650000 ;
      RECT 516.500000 260.350000 549.500000 261.650000 ;
      RECT 507.500000 260.350000 508.500000 261.650000 ;
      RECT 466.500000 260.350000 499.500000 261.650000 ;
      RECT 457.500000 260.350000 458.500000 261.650000 ;
      RECT 416.500000 260.350000 449.500000 261.650000 ;
      RECT 407.500000 260.350000 408.500000 261.650000 ;
      RECT 366.500000 260.350000 399.500000 261.650000 ;
      RECT 357.500000 260.350000 358.500000 261.650000 ;
      RECT 316.500000 260.350000 349.500000 261.650000 ;
      RECT 307.500000 260.350000 308.500000 261.650000 ;
      RECT 266.500000 260.350000 299.500000 261.650000 ;
      RECT 257.500000 260.350000 258.500000 261.650000 ;
      RECT 216.500000 260.350000 249.500000 261.650000 ;
      RECT 207.500000 260.350000 208.500000 261.650000 ;
      RECT 166.500000 260.350000 199.500000 261.650000 ;
      RECT 157.500000 260.350000 158.500000 261.650000 ;
      RECT 116.500000 260.350000 149.500000 261.650000 ;
      RECT 107.500000 260.350000 108.500000 261.650000 ;
      RECT 66.500000 260.350000 99.500000 261.650000 ;
      RECT 57.500000 260.350000 58.500000 261.650000 ;
      RECT 29.500000 260.350000 49.500000 261.650000 ;
      RECT 15.500000 260.350000 16.500000 261.650000 ;
      RECT 0.000000 260.350000 2.500000 263.650000 ;
      RECT 1169.500000 259.650000 1186.000000 260.350000 ;
      RECT 1116.500000 259.650000 1156.500000 260.350000 ;
      RECT 1169.500000 258.350000 1170.500000 259.650000 ;
      RECT 1116.500000 258.350000 1149.500000 259.650000 ;
      RECT 1066.500000 258.350000 1108.500000 260.350000 ;
      RECT 1016.500000 258.350000 1058.500000 260.350000 ;
      RECT 966.500000 258.350000 1008.500000 260.350000 ;
      RECT 916.500000 258.350000 958.500000 260.350000 ;
      RECT 866.500000 258.350000 908.500000 260.350000 ;
      RECT 816.500000 258.350000 858.500000 260.350000 ;
      RECT 766.500000 258.350000 808.500000 260.350000 ;
      RECT 716.500000 258.350000 758.500000 260.350000 ;
      RECT 666.500000 258.350000 708.500000 260.350000 ;
      RECT 616.500000 258.350000 658.500000 260.350000 ;
      RECT 566.500000 258.350000 608.500000 260.350000 ;
      RECT 516.500000 258.350000 558.500000 260.350000 ;
      RECT 466.500000 258.350000 508.500000 260.350000 ;
      RECT 416.500000 258.350000 458.500000 260.350000 ;
      RECT 366.500000 258.350000 408.500000 260.350000 ;
      RECT 316.500000 258.350000 358.500000 260.350000 ;
      RECT 266.500000 258.350000 308.500000 260.350000 ;
      RECT 216.500000 258.350000 258.500000 260.350000 ;
      RECT 166.500000 258.350000 208.500000 260.350000 ;
      RECT 116.500000 258.350000 158.500000 260.350000 ;
      RECT 66.500000 258.350000 108.500000 260.350000 ;
      RECT 29.500000 258.350000 58.500000 260.350000 ;
      RECT 0.000000 258.350000 16.500000 260.350000 ;
      RECT 1157.500000 257.650000 1170.500000 258.350000 ;
      RECT 1183.500000 256.350000 1186.000000 259.650000 ;
      RECT 1169.500000 256.350000 1170.500000 257.650000 ;
      RECT 0.000000 256.350000 1149.500000 258.350000 ;
      RECT 1169.500000 255.650000 1186.000000 256.350000 ;
      RECT 1169.500000 254.350000 1170.500000 255.650000 ;
      RECT 0.000000 254.350000 1156.500000 256.350000 ;
      RECT 0.000000 253.650000 1170.500000 254.350000 ;
      RECT 1183.500000 252.350000 1186.000000 255.650000 ;
      RECT 1169.500000 252.350000 1170.500000 253.650000 ;
      RECT 1169.500000 251.650000 1186.000000 252.350000 ;
      RECT 1169.500000 250.350000 1170.500000 251.650000 ;
      RECT 0.000000 250.350000 1156.500000 253.650000 ;
      RECT 0.000000 249.650000 1170.500000 250.350000 ;
      RECT 1183.500000 248.350000 1186.000000 251.650000 ;
      RECT 1169.500000 248.350000 1170.500000 249.650000 ;
      RECT 1169.500000 247.650000 1186.000000 248.350000 ;
      RECT 1169.500000 246.350000 1170.500000 247.650000 ;
      RECT 0.000000 246.350000 1156.500000 249.650000 ;
      RECT 0.000000 245.650000 1170.500000 246.350000 ;
      RECT 1183.500000 244.350000 1186.000000 247.650000 ;
      RECT 1169.500000 244.350000 1170.500000 245.650000 ;
      RECT 1169.500000 243.650000 1186.000000 244.350000 ;
      RECT 1169.500000 242.350000 1170.500000 243.650000 ;
      RECT 0.000000 242.350000 1156.500000 245.650000 ;
      RECT 0.000000 241.650000 1170.500000 242.350000 ;
      RECT 1183.500000 240.350000 1186.000000 243.650000 ;
      RECT 1169.500000 240.350000 1170.500000 241.650000 ;
      RECT 1169.500000 239.650000 1186.000000 240.350000 ;
      RECT 1169.500000 238.350000 1170.500000 239.650000 ;
      RECT 0.000000 238.350000 1156.500000 241.650000 ;
      RECT 0.000000 237.650000 1170.500000 238.350000 ;
      RECT 1183.500000 236.350000 1186.000000 239.650000 ;
      RECT 1169.500000 236.350000 1170.500000 237.650000 ;
      RECT 1169.500000 235.650000 1186.000000 236.350000 ;
      RECT 1169.500000 234.350000 1170.500000 235.650000 ;
      RECT 0.000000 234.350000 1156.500000 237.650000 ;
      RECT 0.000000 233.650000 1170.500000 234.350000 ;
      RECT 1183.500000 232.350000 1186.000000 235.650000 ;
      RECT 1169.500000 232.350000 1170.500000 233.650000 ;
      RECT 1169.500000 231.650000 1186.000000 232.350000 ;
      RECT 1169.500000 230.350000 1170.500000 231.650000 ;
      RECT 0.000000 230.350000 1156.500000 233.650000 ;
      RECT 0.000000 229.650000 1170.500000 230.350000 ;
      RECT 1183.500000 228.350000 1186.000000 231.650000 ;
      RECT 1169.500000 228.350000 1170.500000 229.650000 ;
      RECT 1169.500000 227.650000 1186.000000 228.350000 ;
      RECT 1169.500000 226.350000 1170.500000 227.650000 ;
      RECT 0.000000 226.350000 1156.500000 229.650000 ;
      RECT 0.000000 225.650000 1170.500000 226.350000 ;
      RECT 1183.500000 224.350000 1186.000000 227.650000 ;
      RECT 1169.500000 224.350000 1170.500000 225.650000 ;
      RECT 1169.500000 223.650000 1186.000000 224.350000 ;
      RECT 1169.500000 222.350000 1170.500000 223.650000 ;
      RECT 0.000000 222.350000 1156.500000 225.650000 ;
      RECT 0.000000 221.650000 1170.500000 222.350000 ;
      RECT 1183.500000 220.350000 1186.000000 223.650000 ;
      RECT 1169.500000 220.350000 1170.500000 221.650000 ;
      RECT 1169.500000 219.650000 1186.000000 220.350000 ;
      RECT 1169.500000 218.350000 1170.500000 219.650000 ;
      RECT 0.000000 218.350000 1156.500000 221.650000 ;
      RECT 0.000000 217.650000 1170.500000 218.350000 ;
      RECT 1183.500000 216.350000 1186.000000 219.650000 ;
      RECT 1169.500000 216.350000 1170.500000 217.650000 ;
      RECT 1169.500000 215.650000 1186.000000 216.350000 ;
      RECT 1169.500000 214.350000 1170.500000 215.650000 ;
      RECT 0.000000 214.350000 1156.500000 217.650000 ;
      RECT 0.000000 213.650000 1170.500000 214.350000 ;
      RECT 1183.500000 212.350000 1186.000000 215.650000 ;
      RECT 1169.500000 212.350000 1170.500000 213.650000 ;
      RECT 1169.500000 211.650000 1186.000000 212.350000 ;
      RECT 1169.500000 210.350000 1170.500000 211.650000 ;
      RECT 0.000000 210.350000 1156.500000 213.650000 ;
      RECT 0.000000 209.650000 1170.500000 210.350000 ;
      RECT 1183.500000 208.350000 1186.000000 211.650000 ;
      RECT 1169.500000 208.350000 1170.500000 209.650000 ;
      RECT 1169.500000 207.650000 1186.000000 208.350000 ;
      RECT 1169.500000 206.350000 1170.500000 207.650000 ;
      RECT 0.000000 206.350000 1156.500000 209.650000 ;
      RECT 0.000000 205.650000 1170.500000 206.350000 ;
      RECT 1183.500000 204.350000 1186.000000 207.650000 ;
      RECT 1169.500000 204.350000 1170.500000 205.650000 ;
      RECT 1169.500000 203.650000 1186.000000 204.350000 ;
      RECT 1169.500000 202.350000 1170.500000 203.650000 ;
      RECT 0.000000 202.350000 1156.500000 205.650000 ;
      RECT 0.000000 201.650000 1170.500000 202.350000 ;
      RECT 1183.500000 200.350000 1186.000000 203.650000 ;
      RECT 1169.500000 200.350000 1170.500000 201.650000 ;
      RECT 1169.500000 199.650000 1186.000000 200.350000 ;
      RECT 1169.500000 198.350000 1170.500000 199.650000 ;
      RECT 0.000000 198.350000 1156.500000 201.650000 ;
      RECT 0.000000 197.650000 1170.500000 198.350000 ;
      RECT 1183.500000 196.350000 1186.000000 199.650000 ;
      RECT 1169.500000 196.350000 1170.500000 197.650000 ;
      RECT 1169.500000 195.650000 1186.000000 196.350000 ;
      RECT 1169.500000 194.350000 1170.500000 195.650000 ;
      RECT 0.000000 194.350000 1156.500000 197.650000 ;
      RECT 0.000000 193.650000 1170.500000 194.350000 ;
      RECT 1183.500000 192.350000 1186.000000 195.650000 ;
      RECT 1169.500000 192.350000 1170.500000 193.650000 ;
      RECT 1169.500000 191.650000 1186.000000 192.350000 ;
      RECT 1169.500000 190.350000 1170.500000 191.650000 ;
      RECT 0.000000 190.350000 1156.500000 193.650000 ;
      RECT 0.000000 189.650000 1170.500000 190.350000 ;
      RECT 1183.500000 188.350000 1186.000000 191.650000 ;
      RECT 1169.500000 188.350000 1170.500000 189.650000 ;
      RECT 1169.500000 187.650000 1186.000000 188.350000 ;
      RECT 1169.500000 186.350000 1170.500000 187.650000 ;
      RECT 0.000000 186.350000 1156.500000 189.650000 ;
      RECT 0.000000 185.650000 1170.500000 186.350000 ;
      RECT 1183.500000 184.350000 1186.000000 187.650000 ;
      RECT 1169.500000 184.350000 1170.500000 185.650000 ;
      RECT 1169.500000 183.650000 1186.000000 184.350000 ;
      RECT 1169.500000 182.350000 1170.500000 183.650000 ;
      RECT 0.000000 182.350000 1156.500000 185.650000 ;
      RECT 0.000000 181.650000 1170.500000 182.350000 ;
      RECT 1183.500000 180.350000 1186.000000 183.650000 ;
      RECT 1169.500000 180.350000 1170.500000 181.650000 ;
      RECT 1169.500000 179.650000 1186.000000 180.350000 ;
      RECT 1169.500000 178.350000 1170.500000 179.650000 ;
      RECT 0.000000 178.350000 1156.500000 181.650000 ;
      RECT 0.000000 177.650000 1170.500000 178.350000 ;
      RECT 1183.500000 176.350000 1186.000000 179.650000 ;
      RECT 1169.500000 176.350000 1170.500000 177.650000 ;
      RECT 1169.500000 175.650000 1186.000000 176.350000 ;
      RECT 1169.500000 174.350000 1170.500000 175.650000 ;
      RECT 0.000000 174.350000 1156.500000 177.650000 ;
      RECT 0.000000 173.650000 1170.500000 174.350000 ;
      RECT 1183.500000 172.350000 1186.000000 175.650000 ;
      RECT 1169.500000 172.350000 1170.500000 173.650000 ;
      RECT 1169.500000 171.650000 1186.000000 172.350000 ;
      RECT 1169.500000 170.350000 1170.500000 171.650000 ;
      RECT 0.000000 170.350000 1156.500000 173.650000 ;
      RECT 0.000000 169.650000 1170.500000 170.350000 ;
      RECT 1183.500000 168.350000 1186.000000 171.650000 ;
      RECT 1169.500000 168.350000 1170.500000 169.650000 ;
      RECT 1169.500000 167.650000 1186.000000 168.350000 ;
      RECT 1169.500000 166.350000 1170.500000 167.650000 ;
      RECT 0.000000 166.350000 1156.500000 169.650000 ;
      RECT 0.000000 165.650000 1170.500000 166.350000 ;
      RECT 1183.500000 164.350000 1186.000000 167.650000 ;
      RECT 1169.500000 164.350000 1170.500000 165.650000 ;
      RECT 1169.500000 163.650000 1186.000000 164.350000 ;
      RECT 1169.500000 162.350000 1170.500000 163.650000 ;
      RECT 0.000000 162.350000 1156.500000 165.650000 ;
      RECT 0.000000 161.650000 1170.500000 162.350000 ;
      RECT 1183.500000 160.350000 1186.000000 163.650000 ;
      RECT 1169.500000 160.350000 1170.500000 161.650000 ;
      RECT 1169.500000 159.650000 1186.000000 160.350000 ;
      RECT 1169.500000 158.350000 1170.500000 159.650000 ;
      RECT 0.000000 158.350000 1156.500000 161.650000 ;
      RECT 0.000000 157.650000 1170.500000 158.350000 ;
      RECT 1183.500000 156.350000 1186.000000 159.650000 ;
      RECT 1169.500000 156.350000 1170.500000 157.650000 ;
      RECT 1169.500000 155.650000 1186.000000 156.350000 ;
      RECT 1169.500000 154.350000 1170.500000 155.650000 ;
      RECT 0.000000 154.350000 1156.500000 157.650000 ;
      RECT 0.000000 153.650000 1170.500000 154.350000 ;
      RECT 1183.500000 152.350000 1186.000000 155.650000 ;
      RECT 1169.500000 152.350000 1170.500000 153.650000 ;
      RECT 1169.500000 151.650000 1186.000000 152.350000 ;
      RECT 1169.500000 150.350000 1170.500000 151.650000 ;
      RECT 0.000000 150.350000 1156.500000 153.650000 ;
      RECT 0.000000 149.650000 1170.500000 150.350000 ;
      RECT 1183.500000 148.350000 1186.000000 151.650000 ;
      RECT 1169.500000 148.350000 1170.500000 149.650000 ;
      RECT 1169.500000 147.650000 1186.000000 148.350000 ;
      RECT 1169.500000 146.350000 1170.500000 147.650000 ;
      RECT 0.000000 146.350000 1156.500000 149.650000 ;
      RECT 0.000000 145.650000 1170.500000 146.350000 ;
      RECT 1183.500000 144.350000 1186.000000 147.650000 ;
      RECT 1169.500000 144.350000 1170.500000 145.650000 ;
      RECT 1169.500000 143.650000 1186.000000 144.350000 ;
      RECT 1169.500000 142.350000 1170.500000 143.650000 ;
      RECT 0.000000 142.350000 1156.500000 145.650000 ;
      RECT 0.000000 141.650000 1170.500000 142.350000 ;
      RECT 1183.500000 140.350000 1186.000000 143.650000 ;
      RECT 1169.500000 140.350000 1170.500000 141.650000 ;
      RECT 1169.500000 139.650000 1186.000000 140.350000 ;
      RECT 1169.500000 138.350000 1170.500000 139.650000 ;
      RECT 0.000000 138.350000 1156.500000 141.650000 ;
      RECT 0.000000 137.650000 1170.500000 138.350000 ;
      RECT 1183.500000 136.350000 1186.000000 139.650000 ;
      RECT 1169.500000 136.350000 1170.500000 137.650000 ;
      RECT 1169.500000 135.650000 1186.000000 136.350000 ;
      RECT 0.000000 135.650000 1156.500000 137.650000 ;
      RECT 1169.500000 134.350000 1170.500000 135.650000 ;
      RECT 1157.500000 133.650000 1170.500000 134.350000 ;
      RECT 1183.500000 132.350000 1186.000000 135.650000 ;
      RECT 1169.500000 132.350000 1170.500000 133.650000 ;
      RECT 0.000000 132.350000 1149.500000 135.650000 ;
      RECT 1169.500000 131.650000 1186.000000 132.350000 ;
      RECT 1169.500000 130.350000 1170.500000 131.650000 ;
      RECT 0.000000 130.350000 1156.500000 132.350000 ;
      RECT 0.000000 129.650000 1170.500000 130.350000 ;
      RECT 1183.500000 128.350000 1186.000000 131.650000 ;
      RECT 1169.500000 128.350000 1170.500000 129.650000 ;
      RECT 1169.500000 127.650000 1186.000000 128.350000 ;
      RECT 1169.500000 126.350000 1170.500000 127.650000 ;
      RECT 0.000000 126.350000 1156.500000 129.650000 ;
      RECT 0.000000 125.650000 1170.500000 126.350000 ;
      RECT 1183.500000 124.350000 1186.000000 127.650000 ;
      RECT 1169.500000 124.350000 1170.500000 125.650000 ;
      RECT 1169.500000 123.650000 1186.000000 124.350000 ;
      RECT 1169.500000 122.350000 1170.500000 123.650000 ;
      RECT 0.000000 122.350000 1156.500000 125.650000 ;
      RECT 0.000000 121.650000 1170.500000 122.350000 ;
      RECT 1183.500000 120.350000 1186.000000 123.650000 ;
      RECT 1169.500000 120.350000 1170.500000 121.650000 ;
      RECT 1169.500000 119.650000 1186.000000 120.350000 ;
      RECT 1169.500000 118.350000 1170.500000 119.650000 ;
      RECT 0.000000 118.350000 1156.500000 121.650000 ;
      RECT 0.000000 117.650000 1170.500000 118.350000 ;
      RECT 1183.500000 116.350000 1186.000000 119.650000 ;
      RECT 1169.500000 116.350000 1170.500000 117.650000 ;
      RECT 1169.500000 115.650000 1186.000000 116.350000 ;
      RECT 1169.500000 114.350000 1170.500000 115.650000 ;
      RECT 0.000000 114.350000 1156.500000 117.650000 ;
      RECT 0.000000 113.650000 1170.500000 114.350000 ;
      RECT 1183.500000 112.350000 1186.000000 115.650000 ;
      RECT 1169.500000 112.350000 1170.500000 113.650000 ;
      RECT 1169.500000 111.650000 1186.000000 112.350000 ;
      RECT 1169.500000 110.350000 1170.500000 111.650000 ;
      RECT 0.000000 110.350000 1156.500000 113.650000 ;
      RECT 0.000000 109.650000 1170.500000 110.350000 ;
      RECT 1183.500000 108.350000 1186.000000 111.650000 ;
      RECT 1169.500000 108.350000 1170.500000 109.650000 ;
      RECT 1169.500000 107.650000 1186.000000 108.350000 ;
      RECT 1169.500000 106.350000 1170.500000 107.650000 ;
      RECT 0.000000 106.350000 1156.500000 109.650000 ;
      RECT 0.000000 105.650000 1170.500000 106.350000 ;
      RECT 1183.500000 104.350000 1186.000000 107.650000 ;
      RECT 1169.500000 104.350000 1170.500000 105.650000 ;
      RECT 1169.500000 103.650000 1186.000000 104.350000 ;
      RECT 1169.500000 102.350000 1170.500000 103.650000 ;
      RECT 0.000000 102.350000 1156.500000 105.650000 ;
      RECT 0.000000 101.650000 1170.500000 102.350000 ;
      RECT 1183.500000 100.350000 1186.000000 103.650000 ;
      RECT 1169.500000 100.350000 1170.500000 101.650000 ;
      RECT 1169.500000 99.650000 1186.000000 100.350000 ;
      RECT 1169.500000 98.350000 1170.500000 99.650000 ;
      RECT 0.000000 98.350000 1156.500000 101.650000 ;
      RECT 0.000000 97.650000 1170.500000 98.350000 ;
      RECT 1183.500000 96.350000 1186.000000 99.650000 ;
      RECT 1169.500000 96.350000 1170.500000 97.650000 ;
      RECT 1169.500000 95.650000 1186.000000 96.350000 ;
      RECT 1169.500000 94.350000 1170.500000 95.650000 ;
      RECT 0.000000 94.350000 1156.500000 97.650000 ;
      RECT 0.000000 93.650000 1170.500000 94.350000 ;
      RECT 1183.500000 92.350000 1186.000000 95.650000 ;
      RECT 1169.500000 92.350000 1170.500000 93.650000 ;
      RECT 1169.500000 91.650000 1186.000000 92.350000 ;
      RECT 1169.500000 90.350000 1170.500000 91.650000 ;
      RECT 0.000000 90.350000 1156.500000 93.650000 ;
      RECT 0.000000 89.650000 1170.500000 90.350000 ;
      RECT 1183.500000 88.350000 1186.000000 91.650000 ;
      RECT 1169.500000 88.350000 1170.500000 89.650000 ;
      RECT 1169.500000 87.650000 1186.000000 88.350000 ;
      RECT 1169.500000 86.350000 1170.500000 87.650000 ;
      RECT 0.000000 86.350000 1156.500000 89.650000 ;
      RECT 0.000000 85.650000 1170.500000 86.350000 ;
      RECT 1183.500000 84.350000 1186.000000 87.650000 ;
      RECT 1169.500000 84.350000 1170.500000 85.650000 ;
      RECT 1169.500000 83.650000 1186.000000 84.350000 ;
      RECT 1169.500000 82.350000 1170.500000 83.650000 ;
      RECT 0.000000 82.350000 1156.500000 85.650000 ;
      RECT 0.000000 81.650000 1170.500000 82.350000 ;
      RECT 1183.500000 80.350000 1186.000000 83.650000 ;
      RECT 1169.500000 80.350000 1170.500000 81.650000 ;
      RECT 1169.500000 79.650000 1186.000000 80.350000 ;
      RECT 1169.500000 78.350000 1170.500000 79.650000 ;
      RECT 0.000000 78.350000 1156.500000 81.650000 ;
      RECT 0.000000 77.650000 1170.500000 78.350000 ;
      RECT 1183.500000 76.350000 1186.000000 79.650000 ;
      RECT 1169.500000 76.350000 1170.500000 77.650000 ;
      RECT 1169.500000 75.650000 1186.000000 76.350000 ;
      RECT 1169.500000 74.350000 1170.500000 75.650000 ;
      RECT 0.000000 74.350000 1156.500000 77.650000 ;
      RECT 0.000000 73.650000 1170.500000 74.350000 ;
      RECT 1183.500000 72.350000 1186.000000 75.650000 ;
      RECT 1169.500000 72.350000 1170.500000 73.650000 ;
      RECT 1169.500000 71.650000 1186.000000 72.350000 ;
      RECT 1169.500000 70.350000 1170.500000 71.650000 ;
      RECT 0.000000 70.350000 1156.500000 73.650000 ;
      RECT 0.000000 69.650000 1170.500000 70.350000 ;
      RECT 1183.500000 68.350000 1186.000000 71.650000 ;
      RECT 1169.500000 68.350000 1170.500000 69.650000 ;
      RECT 1169.500000 67.650000 1186.000000 68.350000 ;
      RECT 1169.500000 66.350000 1170.500000 67.650000 ;
      RECT 0.000000 66.350000 1156.500000 69.650000 ;
      RECT 0.000000 65.650000 1170.500000 66.350000 ;
      RECT 1183.500000 64.350000 1186.000000 67.650000 ;
      RECT 1169.500000 64.350000 1170.500000 65.650000 ;
      RECT 1169.500000 63.650000 1186.000000 64.350000 ;
      RECT 1169.500000 62.350000 1170.500000 63.650000 ;
      RECT 0.000000 62.350000 1156.500000 65.650000 ;
      RECT 0.000000 61.650000 1170.500000 62.350000 ;
      RECT 1183.500000 60.350000 1186.000000 63.650000 ;
      RECT 1169.500000 60.350000 1170.500000 61.650000 ;
      RECT 1169.500000 59.650000 1186.000000 60.350000 ;
      RECT 1169.500000 58.350000 1170.500000 59.650000 ;
      RECT 0.000000 58.350000 1156.500000 61.650000 ;
      RECT 0.000000 57.650000 1170.500000 58.350000 ;
      RECT 1183.500000 56.350000 1186.000000 59.650000 ;
      RECT 1169.500000 56.350000 1170.500000 57.650000 ;
      RECT 1169.500000 55.650000 1186.000000 56.350000 ;
      RECT 1169.500000 54.350000 1170.500000 55.650000 ;
      RECT 0.000000 54.350000 1156.500000 57.650000 ;
      RECT 0.000000 53.650000 1170.500000 54.350000 ;
      RECT 1183.500000 52.350000 1186.000000 55.650000 ;
      RECT 1169.500000 52.350000 1170.500000 53.650000 ;
      RECT 1169.500000 51.650000 1186.000000 52.350000 ;
      RECT 1169.500000 50.350000 1170.500000 51.650000 ;
      RECT 0.000000 50.350000 1156.500000 53.650000 ;
      RECT 0.000000 49.650000 1170.500000 50.350000 ;
      RECT 1183.500000 48.350000 1186.000000 51.650000 ;
      RECT 1169.500000 48.350000 1170.500000 49.650000 ;
      RECT 1169.500000 47.650000 1186.000000 48.350000 ;
      RECT 1169.500000 46.350000 1170.500000 47.650000 ;
      RECT 0.000000 46.350000 1156.500000 49.650000 ;
      RECT 0.000000 45.650000 1170.500000 46.350000 ;
      RECT 1183.500000 44.350000 1186.000000 47.650000 ;
      RECT 1169.500000 44.350000 1170.500000 45.650000 ;
      RECT 1169.500000 43.650000 1186.000000 44.350000 ;
      RECT 1169.500000 42.350000 1170.500000 43.650000 ;
      RECT 0.000000 42.350000 1156.500000 45.650000 ;
      RECT 0.000000 41.650000 1170.500000 42.350000 ;
      RECT 1183.500000 40.350000 1186.000000 43.650000 ;
      RECT 1169.500000 40.350000 1170.500000 41.650000 ;
      RECT 1169.500000 39.650000 1186.000000 40.350000 ;
      RECT 1169.500000 38.350000 1170.500000 39.650000 ;
      RECT 0.000000 38.350000 1156.500000 41.650000 ;
      RECT 0.000000 37.650000 1170.500000 38.350000 ;
      RECT 1183.500000 36.350000 1186.000000 39.650000 ;
      RECT 1169.500000 36.350000 1170.500000 37.650000 ;
      RECT 1169.500000 35.650000 1186.000000 36.350000 ;
      RECT 1169.500000 34.350000 1170.500000 35.650000 ;
      RECT 0.000000 34.350000 1156.500000 37.650000 ;
      RECT 0.000000 33.650000 1170.500000 34.350000 ;
      RECT 1183.500000 32.350000 1186.000000 35.650000 ;
      RECT 1169.500000 32.350000 1170.500000 33.650000 ;
      RECT 1169.500000 31.650000 1186.000000 32.350000 ;
      RECT 1169.500000 30.350000 1170.500000 31.650000 ;
      RECT 0.000000 30.350000 1156.500000 33.650000 ;
      RECT 0.000000 29.650000 1170.500000 30.350000 ;
      RECT 1183.500000 28.350000 1186.000000 31.650000 ;
      RECT 1169.500000 28.350000 1170.500000 29.650000 ;
      RECT 1169.500000 27.650000 1186.000000 28.350000 ;
      RECT 1169.500000 26.350000 1170.500000 27.650000 ;
      RECT 0.000000 26.350000 1156.500000 29.650000 ;
      RECT 0.000000 25.650000 1170.500000 26.350000 ;
      RECT 1183.500000 24.350000 1186.000000 27.650000 ;
      RECT 1169.500000 24.350000 1170.500000 25.650000 ;
      RECT 1169.500000 23.650000 1186.000000 24.350000 ;
      RECT 1169.500000 22.350000 1170.500000 23.650000 ;
      RECT 0.000000 22.350000 1156.500000 25.650000 ;
      RECT 0.000000 21.650000 1170.500000 22.350000 ;
      RECT 1183.500000 20.350000 1186.000000 23.650000 ;
      RECT 1169.500000 20.350000 1170.500000 21.650000 ;
      RECT 1169.500000 19.650000 1186.000000 20.350000 ;
      RECT 1169.500000 18.350000 1170.500000 19.650000 ;
      RECT 0.000000 18.350000 1156.500000 21.650000 ;
      RECT 0.000000 17.650000 1170.500000 18.350000 ;
      RECT 1183.500000 16.350000 1186.000000 19.650000 ;
      RECT 1166.500000 16.350000 1170.500000 17.650000 ;
      RECT 1166.500000 15.650000 1186.000000 16.350000 ;
      RECT 1166.500000 14.350000 1170.500000 15.650000 ;
      RECT 0.000000 14.350000 1158.500000 17.650000 ;
      RECT 0.000000 13.650000 1170.500000 14.350000 ;
      RECT 1183.500000 12.350000 1186.000000 15.650000 ;
      RECT 1166.500000 12.350000 1170.500000 13.650000 ;
      RECT 1166.500000 11.650000 1186.000000 12.350000 ;
      RECT 1166.500000 10.350000 1170.500000 11.650000 ;
      RECT 0.000000 10.350000 1158.500000 13.650000 ;
      RECT 0.000000 9.650000 1170.500000 10.350000 ;
      RECT 1183.500000 8.350000 1186.000000 11.650000 ;
      RECT 1166.500000 8.350000 1170.500000 9.650000 ;
      RECT 1166.500000 7.650000 1186.000000 8.350000 ;
      RECT 1116.500000 7.650000 1158.500000 9.650000 ;
      RECT 1066.500000 7.650000 1108.500000 9.650000 ;
      RECT 1016.500000 7.650000 1058.500000 9.650000 ;
      RECT 966.500000 7.650000 1008.500000 9.650000 ;
      RECT 916.500000 7.650000 958.500000 9.650000 ;
      RECT 866.500000 7.650000 908.500000 9.650000 ;
      RECT 816.500000 7.650000 858.500000 9.650000 ;
      RECT 766.500000 7.650000 808.500000 9.650000 ;
      RECT 716.500000 7.650000 758.500000 9.650000 ;
      RECT 666.500000 7.650000 708.500000 9.650000 ;
      RECT 616.500000 7.650000 658.500000 9.650000 ;
      RECT 566.500000 7.650000 608.500000 9.650000 ;
      RECT 516.500000 7.650000 558.500000 9.650000 ;
      RECT 466.500000 7.650000 508.500000 9.650000 ;
      RECT 416.500000 7.650000 458.500000 9.650000 ;
      RECT 366.500000 7.650000 408.500000 9.650000 ;
      RECT 316.500000 7.650000 358.500000 9.650000 ;
      RECT 266.500000 7.650000 308.500000 9.650000 ;
      RECT 216.500000 7.650000 258.500000 9.650000 ;
      RECT 166.500000 7.650000 208.500000 9.650000 ;
      RECT 116.500000 7.650000 158.500000 9.650000 ;
      RECT 66.500000 7.650000 108.500000 9.650000 ;
      RECT 0.000000 7.650000 58.500000 9.650000 ;
      RECT 1166.500000 6.350000 1170.500000 7.650000 ;
      RECT 1157.500000 6.350000 1158.500000 7.650000 ;
      RECT 1116.500000 6.350000 1149.500000 7.650000 ;
      RECT 1107.500000 6.350000 1108.500000 7.650000 ;
      RECT 1066.500000 6.350000 1099.500000 7.650000 ;
      RECT 1057.500000 6.350000 1058.500000 7.650000 ;
      RECT 1016.500000 6.350000 1049.500000 7.650000 ;
      RECT 1007.500000 6.350000 1008.500000 7.650000 ;
      RECT 966.500000 6.350000 999.500000 7.650000 ;
      RECT 957.500000 6.350000 958.500000 7.650000 ;
      RECT 916.500000 6.350000 949.500000 7.650000 ;
      RECT 907.500000 6.350000 908.500000 7.650000 ;
      RECT 866.500000 6.350000 899.500000 7.650000 ;
      RECT 857.500000 6.350000 858.500000 7.650000 ;
      RECT 816.500000 6.350000 849.500000 7.650000 ;
      RECT 807.500000 6.350000 808.500000 7.650000 ;
      RECT 766.500000 6.350000 799.500000 7.650000 ;
      RECT 757.500000 6.350000 758.500000 7.650000 ;
      RECT 716.500000 6.350000 749.500000 7.650000 ;
      RECT 707.500000 6.350000 708.500000 7.650000 ;
      RECT 666.500000 6.350000 699.500000 7.650000 ;
      RECT 657.500000 6.350000 658.500000 7.650000 ;
      RECT 616.500000 6.350000 649.500000 7.650000 ;
      RECT 607.500000 6.350000 608.500000 7.650000 ;
      RECT 566.500000 6.350000 599.500000 7.650000 ;
      RECT 557.500000 6.350000 558.500000 7.650000 ;
      RECT 516.500000 6.350000 549.500000 7.650000 ;
      RECT 507.500000 6.350000 508.500000 7.650000 ;
      RECT 466.500000 6.350000 499.500000 7.650000 ;
      RECT 457.500000 6.350000 458.500000 7.650000 ;
      RECT 416.500000 6.350000 449.500000 7.650000 ;
      RECT 407.500000 6.350000 408.500000 7.650000 ;
      RECT 366.500000 6.350000 399.500000 7.650000 ;
      RECT 357.500000 6.350000 358.500000 7.650000 ;
      RECT 316.500000 6.350000 349.500000 7.650000 ;
      RECT 307.500000 6.350000 308.500000 7.650000 ;
      RECT 266.500000 6.350000 299.500000 7.650000 ;
      RECT 257.500000 6.350000 258.500000 7.650000 ;
      RECT 216.500000 6.350000 249.500000 7.650000 ;
      RECT 207.500000 6.350000 208.500000 7.650000 ;
      RECT 166.500000 6.350000 199.500000 7.650000 ;
      RECT 157.500000 6.350000 158.500000 7.650000 ;
      RECT 116.500000 6.350000 149.500000 7.650000 ;
      RECT 107.500000 6.350000 108.500000 7.650000 ;
      RECT 66.500000 6.350000 99.500000 7.650000 ;
      RECT 57.500000 6.350000 58.500000 7.650000 ;
      RECT 1157.500000 5.650000 1170.500000 6.350000 ;
      RECT 1107.500000 5.650000 1149.500000 6.350000 ;
      RECT 1057.500000 5.650000 1099.500000 6.350000 ;
      RECT 1007.500000 5.650000 1049.500000 6.350000 ;
      RECT 957.500000 5.650000 999.500000 6.350000 ;
      RECT 907.500000 5.650000 949.500000 6.350000 ;
      RECT 857.500000 5.650000 899.500000 6.350000 ;
      RECT 807.500000 5.650000 849.500000 6.350000 ;
      RECT 757.500000 5.650000 799.500000 6.350000 ;
      RECT 707.500000 5.650000 749.500000 6.350000 ;
      RECT 657.500000 5.650000 699.500000 6.350000 ;
      RECT 607.500000 5.650000 649.500000 6.350000 ;
      RECT 557.500000 5.650000 599.500000 6.350000 ;
      RECT 507.500000 5.650000 549.500000 6.350000 ;
      RECT 457.500000 5.650000 499.500000 6.350000 ;
      RECT 407.500000 5.650000 449.500000 6.350000 ;
      RECT 357.500000 5.650000 399.500000 6.350000 ;
      RECT 307.500000 5.650000 349.500000 6.350000 ;
      RECT 257.500000 5.650000 299.500000 6.350000 ;
      RECT 207.500000 5.650000 249.500000 6.350000 ;
      RECT 157.500000 5.650000 199.500000 6.350000 ;
      RECT 107.500000 5.650000 149.500000 6.350000 ;
      RECT 57.500000 5.650000 99.500000 6.350000 ;
      RECT 1183.500000 4.350000 1186.000000 7.650000 ;
      RECT 1166.500000 4.350000 1170.500000 5.650000 ;
      RECT 1157.500000 4.350000 1158.500000 5.650000 ;
      RECT 1116.500000 4.350000 1149.500000 5.650000 ;
      RECT 1107.500000 4.350000 1108.500000 5.650000 ;
      RECT 1066.500000 4.350000 1099.500000 5.650000 ;
      RECT 1057.500000 4.350000 1058.500000 5.650000 ;
      RECT 1016.500000 4.350000 1049.500000 5.650000 ;
      RECT 1007.500000 4.350000 1008.500000 5.650000 ;
      RECT 966.500000 4.350000 999.500000 5.650000 ;
      RECT 957.500000 4.350000 958.500000 5.650000 ;
      RECT 916.500000 4.350000 949.500000 5.650000 ;
      RECT 907.500000 4.350000 908.500000 5.650000 ;
      RECT 866.500000 4.350000 899.500000 5.650000 ;
      RECT 857.500000 4.350000 858.500000 5.650000 ;
      RECT 816.500000 4.350000 849.500000 5.650000 ;
      RECT 807.500000 4.350000 808.500000 5.650000 ;
      RECT 766.500000 4.350000 799.500000 5.650000 ;
      RECT 757.500000 4.350000 758.500000 5.650000 ;
      RECT 716.500000 4.350000 749.500000 5.650000 ;
      RECT 707.500000 4.350000 708.500000 5.650000 ;
      RECT 666.500000 4.350000 699.500000 5.650000 ;
      RECT 657.500000 4.350000 658.500000 5.650000 ;
      RECT 616.500000 4.350000 649.500000 5.650000 ;
      RECT 607.500000 4.350000 608.500000 5.650000 ;
      RECT 566.500000 4.350000 599.500000 5.650000 ;
      RECT 557.500000 4.350000 558.500000 5.650000 ;
      RECT 516.500000 4.350000 549.500000 5.650000 ;
      RECT 507.500000 4.350000 508.500000 5.650000 ;
      RECT 466.500000 4.350000 499.500000 5.650000 ;
      RECT 457.500000 4.350000 458.500000 5.650000 ;
      RECT 416.500000 4.350000 449.500000 5.650000 ;
      RECT 407.500000 4.350000 408.500000 5.650000 ;
      RECT 366.500000 4.350000 399.500000 5.650000 ;
      RECT 357.500000 4.350000 358.500000 5.650000 ;
      RECT 316.500000 4.350000 349.500000 5.650000 ;
      RECT 307.500000 4.350000 308.500000 5.650000 ;
      RECT 266.500000 4.350000 299.500000 5.650000 ;
      RECT 257.500000 4.350000 258.500000 5.650000 ;
      RECT 216.500000 4.350000 249.500000 5.650000 ;
      RECT 207.500000 4.350000 208.500000 5.650000 ;
      RECT 166.500000 4.350000 199.500000 5.650000 ;
      RECT 157.500000 4.350000 158.500000 5.650000 ;
      RECT 116.500000 4.350000 149.500000 5.650000 ;
      RECT 107.500000 4.350000 108.500000 5.650000 ;
      RECT 66.500000 4.350000 99.500000 5.650000 ;
      RECT 57.500000 4.350000 58.500000 5.650000 ;
      RECT 15.500000 4.350000 49.500000 7.650000 ;
      RECT 0.000000 4.350000 2.500000 7.650000 ;
      RECT 1116.500000 3.650000 1158.500000 4.350000 ;
      RECT 1066.500000 3.650000 1108.500000 4.350000 ;
      RECT 1016.500000 3.650000 1058.500000 4.350000 ;
      RECT 966.500000 3.650000 1008.500000 4.350000 ;
      RECT 916.500000 3.650000 958.500000 4.350000 ;
      RECT 866.500000 3.650000 908.500000 4.350000 ;
      RECT 816.500000 3.650000 858.500000 4.350000 ;
      RECT 766.500000 3.650000 808.500000 4.350000 ;
      RECT 716.500000 3.650000 758.500000 4.350000 ;
      RECT 666.500000 3.650000 708.500000 4.350000 ;
      RECT 616.500000 3.650000 658.500000 4.350000 ;
      RECT 566.500000 3.650000 608.500000 4.350000 ;
      RECT 516.500000 3.650000 558.500000 4.350000 ;
      RECT 466.500000 3.650000 508.500000 4.350000 ;
      RECT 416.500000 3.650000 458.500000 4.350000 ;
      RECT 366.500000 3.650000 408.500000 4.350000 ;
      RECT 316.500000 3.650000 358.500000 4.350000 ;
      RECT 266.500000 3.650000 308.500000 4.350000 ;
      RECT 216.500000 3.650000 258.500000 4.350000 ;
      RECT 166.500000 3.650000 208.500000 4.350000 ;
      RECT 116.500000 3.650000 158.500000 4.350000 ;
      RECT 66.500000 3.650000 108.500000 4.350000 ;
      RECT 0.000000 3.650000 58.500000 4.350000 ;
      RECT 1166.500000 2.350000 1186.000000 4.350000 ;
      RECT 1157.500000 2.350000 1158.500000 3.650000 ;
      RECT 1116.500000 2.350000 1149.500000 3.650000 ;
      RECT 1107.500000 2.350000 1108.500000 3.650000 ;
      RECT 1066.500000 2.350000 1099.500000 3.650000 ;
      RECT 1057.500000 2.350000 1058.500000 3.650000 ;
      RECT 1016.500000 2.350000 1049.500000 3.650000 ;
      RECT 1007.500000 2.350000 1008.500000 3.650000 ;
      RECT 966.500000 2.350000 999.500000 3.650000 ;
      RECT 957.500000 2.350000 958.500000 3.650000 ;
      RECT 916.500000 2.350000 949.500000 3.650000 ;
      RECT 907.500000 2.350000 908.500000 3.650000 ;
      RECT 866.500000 2.350000 899.500000 3.650000 ;
      RECT 857.500000 2.350000 858.500000 3.650000 ;
      RECT 816.500000 2.350000 849.500000 3.650000 ;
      RECT 807.500000 2.350000 808.500000 3.650000 ;
      RECT 766.500000 2.350000 799.500000 3.650000 ;
      RECT 757.500000 2.350000 758.500000 3.650000 ;
      RECT 716.500000 2.350000 749.500000 3.650000 ;
      RECT 707.500000 2.350000 708.500000 3.650000 ;
      RECT 666.500000 2.350000 699.500000 3.650000 ;
      RECT 657.500000 2.350000 658.500000 3.650000 ;
      RECT 616.500000 2.350000 649.500000 3.650000 ;
      RECT 607.500000 2.350000 608.500000 3.650000 ;
      RECT 566.500000 2.350000 599.500000 3.650000 ;
      RECT 557.500000 2.350000 558.500000 3.650000 ;
      RECT 516.500000 2.350000 549.500000 3.650000 ;
      RECT 507.500000 2.350000 508.500000 3.650000 ;
      RECT 466.500000 2.350000 499.500000 3.650000 ;
      RECT 457.500000 2.350000 458.500000 3.650000 ;
      RECT 416.500000 2.350000 449.500000 3.650000 ;
      RECT 407.500000 2.350000 408.500000 3.650000 ;
      RECT 366.500000 2.350000 399.500000 3.650000 ;
      RECT 357.500000 2.350000 358.500000 3.650000 ;
      RECT 316.500000 2.350000 349.500000 3.650000 ;
      RECT 307.500000 2.350000 308.500000 3.650000 ;
      RECT 266.500000 2.350000 299.500000 3.650000 ;
      RECT 257.500000 2.350000 258.500000 3.650000 ;
      RECT 216.500000 2.350000 249.500000 3.650000 ;
      RECT 207.500000 2.350000 208.500000 3.650000 ;
      RECT 166.500000 2.350000 199.500000 3.650000 ;
      RECT 157.500000 2.350000 158.500000 3.650000 ;
      RECT 116.500000 2.350000 149.500000 3.650000 ;
      RECT 107.500000 2.350000 108.500000 3.650000 ;
      RECT 66.500000 2.350000 99.500000 3.650000 ;
      RECT 57.500000 2.350000 58.500000 3.650000 ;
      RECT 1157.500000 0.350000 1186.000000 2.350000 ;
      RECT 1107.500000 0.350000 1149.500000 2.350000 ;
      RECT 1057.500000 0.350000 1099.500000 2.350000 ;
      RECT 1007.500000 0.350000 1049.500000 2.350000 ;
      RECT 957.500000 0.350000 999.500000 2.350000 ;
      RECT 907.500000 0.350000 949.500000 2.350000 ;
      RECT 857.500000 0.350000 899.500000 2.350000 ;
      RECT 807.500000 0.350000 849.500000 2.350000 ;
      RECT 757.500000 0.350000 799.500000 2.350000 ;
      RECT 707.500000 0.350000 749.500000 2.350000 ;
      RECT 657.500000 0.350000 699.500000 2.350000 ;
      RECT 607.500000 0.350000 649.500000 2.350000 ;
      RECT 557.500000 0.350000 599.500000 2.350000 ;
      RECT 507.500000 0.350000 549.500000 2.350000 ;
      RECT 457.500000 0.350000 499.500000 2.350000 ;
      RECT 407.500000 0.350000 449.500000 2.350000 ;
      RECT 357.500000 0.350000 399.500000 2.350000 ;
      RECT 307.500000 0.350000 349.500000 2.350000 ;
      RECT 257.500000 0.350000 299.500000 2.350000 ;
      RECT 207.500000 0.350000 249.500000 2.350000 ;
      RECT 157.500000 0.350000 199.500000 2.350000 ;
      RECT 107.500000 0.350000 149.500000 2.350000 ;
      RECT 57.500000 0.350000 99.500000 2.350000 ;
      RECT 0.000000 0.350000 49.500000 3.650000 ;
      RECT 0.000000 0.000000 1186.000000 0.350000 ;
  END
END MCU

END LIBRARY
