/home/mseminario2/chips/myshkin/ip/rom_hvt_pg/rom_hvt_pg.lef