

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO MCU 
  PIN resetn_in 
    ANTENNAPARTIALMETALAREA 0.9625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.235 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.658 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9392 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 24.822 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 109.261 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 939.327 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4139.7 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6 ;
  END resetn_in
  PIN resetn_out 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.301 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3684 LAYER M2 ;
  END resetn_out
  PIN resetn_dir 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6654 LAYER M2 ;
  END resetn_dir
  PIN resetn_ren 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6378 LAYER M2 ;
  END resetn_ren
  PIN prt1_in[7] 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.464 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.7296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 207.026 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 887.026 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt1_in[7]
  PIN prt1_in[6] 
    ANTENNAPARTIALMETALAREA 1.3925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.127 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.588 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.4752 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 468.035 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2062.77 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3 ;
  END prt1_in[6]
  PIN prt1_in[5] 
    ANTENNAPARTIALMETALAREA 1.0325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.543 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.548 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.2992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 323.159 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1414.36 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END prt1_in[5]
  PIN prt1_in[4] 
    ANTENNAPARTIALMETALAREA 6.1125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.895 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.646 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.0864 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3232 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2577 LAYER M4 ; 
    ANTENNAMAXAREACAR 14.4498 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 63.3398 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.943396 LAYER VIA4 ;
  END prt1_in[4]
  PIN prt1_in[3] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.016 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.8742 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.9686 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.628931 LAYER VIA3 ;
  END prt1_in[3]
  PIN prt1_in[2] 
    ANTENNAPARTIALMETALAREA 4.5975 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.273 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 14.448 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.6592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1449 LAYER M3 ; 
    ANTENNAMAXAREACAR 123.243 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 541.326 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.956084 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.422 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3008 LAYER M4 ;
    ANTENNAGATEAREA 0.2118 LAYER M4 ; 
    ANTENNAMAXAREACAR 129.957 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 571.075 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.956084 LAYER VIA4 ;
  END prt1_in[2]
  PIN prt1_in[1] 
    ANTENNAPARTIALMETALAREA 13.1935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.0954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.926 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.9184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0481 LAYER M3 ; 
    ANTENNAMAXAREACAR 272.119 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1197.84 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.831601 LAYER VIA3 ;
  END prt1_in[1]
  PIN prt1_in[0] 
    ANTENNAPARTIALMETALAREA 17.3555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 76.3642 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0447 LAYER M2 ; 
    ANTENNAMAXAREACAR 451.109 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 1959.53 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.447427 LAYER VIA2 ;
  END prt1_in[0]
  PIN prt1_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.414 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.4656 LAYER M2 ;
  END prt1_out[7]
  PIN prt1_out[6] 
    ANTENNAPARTIALMETALAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5584 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.198 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9152 LAYER M3 ;
  END prt1_out[6]
  PIN prt1_out[5] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[5]
  PIN prt1_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[4]
  PIN prt1_out[3] 
    ANTENNAPARTIALMETALAREA 0.976 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2944 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.982 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.9648 LAYER M3 ;
  END prt1_out[3]
  PIN prt1_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[2]
  PIN prt1_out[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END prt1_out[1]
  PIN prt1_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.175 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.258 LAYER M2 ;
  END prt1_out[0]
  PIN prt1_dir[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[7]
  PIN prt1_dir[6] 
    ANTENNAPARTIALMETALAREA 0.3565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5686 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4784 LAYER M3 ;
  END prt1_dir[6]
  PIN prt1_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
  END prt1_dir[5]
  PIN prt1_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
  END prt1_dir[4]
  PIN prt1_dir[3] 
    ANTENNAPARTIALMETALAREA 0.7165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1526 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.966 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.8944 LAYER M3 ;
  END prt1_dir[3]
  PIN prt1_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6842 LAYER M2 ;
  END prt1_dir[2]
  PIN prt1_dir[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[1]
  PIN prt1_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.4745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.5758 LAYER M2 ;
  END prt1_dir[0]
  PIN prt1_ren[7] 
    ANTENNAPARTIALMETALAREA 0.0805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3542 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.486 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5824 LAYER M3 ;
  END prt1_ren[7]
  PIN prt1_ren[6] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.146 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M3 ;
  END prt1_ren[6]
  PIN prt1_ren[5] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
  END prt1_ren[5]
  PIN prt1_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2 ;
  END prt1_ren[4]
  PIN prt1_ren[3] 
    ANTENNAPARTIALMETALAREA 0.2475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.089 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.902 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.0128 LAYER M3 ;
  END prt1_ren[3]
  PIN prt1_ren[2] 
    ANTENNAPARTIALMETALAREA 3.6935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.2954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.626 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9984 LAYER M3 ;
  END prt1_ren[2]
  PIN prt1_ren[1] 
    ANTENNAPARTIALMETALAREA 8.3915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.9226 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.484 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.038 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6112 LAYER M4 ;
  END prt1_ren[1]
  PIN prt1_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.9505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 52.6702 LAYER M2 ;
  END prt1_ren[0]
  PIN prt2_in[7] 
    ANTENNAPARTIALMETALAREA 0.8145 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6278 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0595 LAYER M2 ; 
    ANTENNAMAXAREACAR 14.6437 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 64.3597 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.336134 LAYER VIA2 ;
  END prt2_in[7]
  PIN prt2_in[6] 
    ANTENNAPARTIALMETALAREA 0.7005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1262 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 23.098 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 100.83 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END prt2_in[6]
  PIN prt2_in[5] 
    ANTENNAPARTIALMETALAREA 0.2785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2254 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 LAYER M2 ; 
    ANTENNAMAXAREACAR 4.20556 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 17.2796 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.185185 LAYER VIA2 ;
  END prt2_in[5]
  PIN prt2_in[4] 
    ANTENNAPARTIALMETALAREA 0.8445 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7598 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 7.2728 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 31.6242 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2 ;
  END prt2_in[4]
  PIN prt2_in[3] 
    ANTENNAPARTIALMETALAREA 0.174 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1914 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.244 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4444 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 3.04 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.696 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M4 ; 
    ANTENNAMAXAREACAR 27.3487 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 37.6462 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.471698 LAYER VIA4 ;
  END prt2_in[3]
  PIN prt2_in[2] 
    ANTENNAPARTIALMETALAREA 0.7155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1482 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0893 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.37514 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 40.0112 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.223964 LAYER VIA2 ;
  END prt2_in[2]
  PIN prt2_in[1] 
    ANTENNAPARTIALMETALAREA 0.4555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0042 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0671 LAYER M2 ; 
    ANTENNAMAXAREACAR 8.26006 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 35.2876 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.298063 LAYER VIA2 ;
  END prt2_in[1]
  PIN prt2_in[0] 
    ANTENNAPARTIALMETALAREA 0.5335 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3914 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M2 ; 
    ANTENNAMAXAREACAR 4.89413 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 20.5996 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.104822 LAYER VIA2 ;
  END prt2_in[0]
  PIN prt2_out[7] 
    ANTENNAPARTIALMETALAREA 0.631 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0368 LAYER M3 ;
  END prt2_out[7]
  PIN prt2_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.717 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1988 LAYER M2 ;
  END prt2_out[6]
  PIN prt2_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.579 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6356 LAYER M2 ;
  END prt2_out[5]
  PIN prt2_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.297 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3508 LAYER M2 ;
  END prt2_out[4]
  PIN prt2_out[3] 
    ANTENNAPARTIALMETALAREA 0.452 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.126 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.1984 LAYER M3 ;
  END prt2_out[3]
  PIN prt2_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2 ;
  END prt2_out[2]
  PIN prt2_out[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.279 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2276 LAYER M2 ;
  END prt2_out[1]
  PIN prt2_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.512 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M2 ;
  END prt2_out[0]
  PIN prt2_dir[7] 
    ANTENNAPARTIALMETALAREA 0.691 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.002 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6528 LAYER M3 ;
  END prt2_dir[7]
  PIN prt2_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6334 LAYER M2 ;
  END prt2_dir[6]
  PIN prt2_dir[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1198 LAYER M2 ;
  END prt2_dir[5]
  PIN prt2_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3486 LAYER M2 ;
  END prt2_dir[4]
  PIN prt2_dir[3] 
    ANTENNAPARTIALMETALAREA 0.3315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4586 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.446 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.6064 LAYER M3 ;
  END prt2_dir[3]
  PIN prt2_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3706 LAYER M2 ;
  END prt2_dir[2]
  PIN prt2_dir[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0778 LAYER M2 ;
  END prt2_dir[1]
  PIN prt2_dir[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3882 LAYER M2 ;
  END prt2_dir[0]
  PIN prt2_ren[7] 
    ANTENNAPARTIALMETALAREA 0.7435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2714 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9008 LAYER M3 ;
  END prt2_ren[7]
  PIN prt2_ren[6] 
    ANTENNAPARTIALMETALAREA 0.5945 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6158 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
  END prt2_ren[6]
  PIN prt2_ren[5] 
    ANTENNAPARTIALMETALAREA 0.6105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6862 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.962 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.4768 LAYER M3 ;
  END prt2_ren[5]
  PIN prt2_ren[4] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3034 LAYER M2 ;
  END prt2_ren[4]
  PIN prt2_ren[3] 
    ANTENNAPARTIALMETALAREA 0.5505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.2528 LAYER M3 ;
  END prt2_ren[3]
  PIN prt2_ren[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2078 LAYER M2 ;
  END prt2_ren[2]
  PIN prt2_ren[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.243 LAYER M2 ;
  END prt2_ren[1]
  PIN prt2_ren[0] 
    ANTENNAPARTIALMETALAREA 0.3675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.9328 LAYER M3 ;
  END prt2_ren[0]
  PIN prt3_in[7] 
    ANTENNAPARTIALMETALAREA 24.7525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 108.911 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.606 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.5104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 504.945 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2208.71 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[7]
  PIN prt3_in[6] 
    ANTENNAPARTIALMETALAREA 15.8905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 69.9622 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 587.98 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2587.28 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2 ;
  END prt3_in[6]
  PIN prt3_in[5] 
    ANTENNAPARTIALMETALAREA 6.8165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.9926 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.484 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.604 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5456 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 396.469 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1747.23 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.89702 LAYER VIA4 ;
  END prt3_in[5]
  PIN prt3_in[4] 
    ANTENNAPARTIALMETALAREA 0.4925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.167 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.6848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 144.627 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 634.569 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.734684 LAYER VIA3 ;
  END prt3_in[4]
  PIN prt3_in[3] 
    ANTENNAPARTIALMETALAREA 3.8935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.4048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 LAYER M3 ; 
    ANTENNAMAXAREACAR 112.461 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 493.461 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.734684 LAYER VIA3 ;
  END prt3_in[3]
  PIN prt3_in[2] 
    ANTENNAPARTIALMETALAREA 10.9355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 48.2042 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.484 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0752 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M4 ; 
    ANTENNAMAXAREACAR 68.7731 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 306.015 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.84502 LAYER VIA4 ;
  END prt3_in[2]
  PIN prt3_in[1] 
    ANTENNAPARTIALMETALAREA 22.8695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 100.758 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M2 ; 
    ANTENNAMAXAREACAR 621.016 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2735.59 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.186 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M3 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 622.808 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2743.9 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3 ;
  END prt3_in[1]
  PIN prt3_in[0] 
    ANTENNAPARTIALMETALAREA 1.8745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2918 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.498 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.8352 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 296.87 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1290.32 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt3_in[0]
  PIN prt3_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.975 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 66.066 LAYER M2 ;
  END prt3_out[7]
  PIN prt3_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.983 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.4132 LAYER M2 ;
  END prt3_out[6]
  PIN prt3_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.241 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1044 LAYER M2 ;
  END prt3_out[5]
  PIN prt3_out[4] 
    ANTENNAPARTIALMETALAREA 1.938 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5712 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.9568 LAYER M3 ;
  END prt3_out[4]
  PIN prt3_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3124 LAYER M2 ;
  END prt3_out[3]
  PIN prt3_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 8.019 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.3716 LAYER M2 ;
  END prt3_out[2]
  PIN prt3_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.999 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 57.2836 LAYER M2 ;
  END prt3_out[1]
  PIN prt3_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.041 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.8244 LAYER M2 ;
  END prt3_out[0]
  PIN prt3_dir[7] 
    ANTENNAPARTIALMETALAREA 13.8765 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.0566 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3968 LAYER M3 ;
  END prt3_dir[7]
  PIN prt3_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.9498 LAYER M2 ;
  END prt3_dir[6]
  PIN prt3_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt3_dir[5]
  PIN prt3_dir[4] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
  END prt3_dir[4]
  PIN prt3_dir[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt3_dir[3]
  PIN prt3_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.1165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6446 LAYER M2 ;
  END prt3_dir[2]
  PIN prt3_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.9965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.6286 LAYER M2 ;
  END prt3_dir[1]
  PIN prt3_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.0435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.4794 LAYER M2 ;
  END prt3_dir[0]
  PIN prt3_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.4035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.0634 LAYER M2 ;
  END prt3_ren[7]
  PIN prt3_ren[6] 
    ANTENNAPARTIALMETALAREA 0.5805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5542 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.816 LAYER M3 ;
  END prt3_ren[6]
  PIN prt3_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.4615 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5626 LAYER M2 ;
  END prt3_ren[5]
  PIN prt3_ren[4] 
    ANTENNAPARTIALMETALAREA 0.2605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1462 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.138 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2512 LAYER M3 ;
  END prt3_ren[4]
  PIN prt3_ren[3] 
    ANTENNAPARTIALMETALAREA 0.0475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.209 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.984 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.6176 LAYER M3 ;
  END prt3_ren[3]
  PIN prt3_ren[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 9.6505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 42.5502 LAYER M2 ;
  END prt3_ren[2]
  PIN prt3_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.3925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 63.459 LAYER M2 ;
  END prt3_ren[1]
  PIN prt3_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.5255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2442 LAYER M2 ;
  END prt3_ren[0]
  PIN prt4_in[7] 
    ANTENNAPARTIALMETALAREA 2.8755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6522 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 27.896 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 122.918 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1456 LAYER M3 ; 
    ANTENNAMAXAREACAR 204.646 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 900.794 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
  END prt4_in[7]
  PIN prt4_in[6] 
    ANTENNAPARTIALMETALAREA 1.6355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1962 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 17.944 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 79.0416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 284.081 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1248.19 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
  END prt4_in[6]
  PIN prt4_in[5] 
    ANTENNAPARTIALMETALAREA 2.3155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.528 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.0112 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 110.891 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 482.45 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.27669 LAYER VIA3 ;
  END prt4_in[5]
  PIN prt4_in[4] 
    ANTENNAPARTIALMETALAREA 4.3355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0762 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.145 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 120.358 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9632 LAYER M4 ;
    ANTENNAGATEAREA 0.1204 LAYER M4 ; 
    ANTENNAMAXAREACAR 36.4307 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 161.58 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA4 ;
  END prt4_in[4]
  PIN prt4_in[3] 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.418 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.0832 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 5.678 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.0272 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1456 LAYER M4 ; 
    ANTENNAMAXAREACAR 48.2889 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 212.608 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.22137 LAYER VIA4 ;
  END prt4_in[3]
  PIN prt4_in[2] 
    ANTENNAPARTIALMETALAREA 5.8925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.015 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M2 ; 
    ANTENNAMAXAREACAR 61.6906 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 270.041 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.542005 LAYER VIA2 ;
  END prt4_in[2]
  PIN prt4_in[1] 
    ANTENNAPARTIALMETALAREA 0.731 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 20.778 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.4672 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 7.598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.4752 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 87.8771 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 387.104 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA4 ;
  END prt4_in[1]
  PIN prt4_in[0] 
    ANTENNAPARTIALMETALAREA 0.2725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 27.886 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 122.742 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 1077.86 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4725.82 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt4_in[0]
  PIN prt4_out[7] 
    ANTENNAPARTIALMETALAREA 10.092 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1606 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 46.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.48 LAYER M3 ;
  END prt4_out[7]
  PIN prt4_out[6] 
    ANTENNAPARTIALMETALAREA 8.492 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4006 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 32.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.728 LAYER M3 ;
  END prt4_out[6]
  PIN prt4_out[5] 
    ANTENNAPARTIALMETALAREA 0.43 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.473 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 19.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.088 LAYER M3 ;
  END prt4_out[5]
  PIN prt4_out[4] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.8902 LAYER M3 ;
  END prt4_out[4]
  PIN prt4_out[3] 
    ANTENNAPARTIALMETALAREA 0.939 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1316 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.806 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.5904 LAYER M3 ;
  END prt4_out[3]
  PIN prt4_out[2] 
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.0608 LAYER M3 ;
  END prt4_out[2]
  PIN prt4_out[1] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.962 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 74.6768 LAYER M6 ;
  END prt4_out[1]
  PIN prt4_out[0] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[0]
  PIN prt4_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4366 LAYER M2 ;
  END prt4_dir[7]
  PIN prt4_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2286 LAYER M2 ;
  END prt4_dir[6]
  PIN prt4_dir[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3222 LAYER M2 ;
  END prt4_dir[5]
  PIN prt4_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3814 LAYER M2 ;
  END prt4_dir[4]
  PIN prt4_dir[3] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7008 LAYER M3 ;
  END prt4_dir[3]
  PIN prt4_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.6395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3018 LAYER M2 ;
  END prt4_dir[2]
  PIN prt4_dir[1] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.722 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.6208 LAYER M6 ;
  END prt4_dir[1]
  PIN prt4_dir[0] 
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.962 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.2768 LAYER M6 ;
  END prt4_dir[0]
  PIN prt4_ren[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3178 LAYER M2 ;
  END prt4_ren[7]
  PIN prt4_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.497 LAYER M2 ;
  END prt4_ren[6]
  PIN prt4_ren[5] 
    ANTENNAPARTIALMETALAREA 0.6505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8622 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.766 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.2144 LAYER M3 ;
  END prt4_ren[5]
  PIN prt4_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.6825 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.447 LAYER M2 ;
  END prt4_ren[4]
  PIN prt4_ren[3] 
    ANTENNAPARTIALMETALAREA 0.9035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.142 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2688 LAYER M3 ;
  END prt4_ren[3]
  PIN prt4_ren[2] 
    ANTENNAPARTIALMETALAREA 0.6635 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9194 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.4608 LAYER M3 ;
  END prt4_ren[2]
  PIN prt4_ren[1] 
    ANTENNAPARTIALMETALAREA 0.8035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6 ;
  END prt4_ren[1]
  PIN prt4_ren[0] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 17.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 75.3808 LAYER M6 ;
  END prt4_ren[0]
  PIN use_dac_glb_bias 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3222 LAYER M2 ;
  END use_dac_glb_bias
  PIN en_bias_buf 
    ANTENNAPARTIALMETALAREA 0.076 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.998 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 26.4352 LAYER M6 ;
  END en_bias_buf
  PIN en_bias_gen 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.429 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9316 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.926 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.3184 LAYER M6 ;
  END en_bias_gen
  PIN BIAS_ADJ[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4 LAYER M3 ;
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.728 LAYER M3 ;
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.162 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M4 ;
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2] 
    ANTENNAPARTIALMETALAREA 2.07 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.152 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.918 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0832 LAYER M3 ;
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0645 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3278 LAYER M2 ;
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.584 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8576 LAYER M2 ;
  END BIAS_DBP[13]
  PIN BIAS_DBP[12] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.098 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8752 LAYER M5 ;
  END BIAS_DBP[12]
  PIN BIAS_DBP[11] 
    ANTENNAPARTIALMETALAREA 0.05 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.428 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9712 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.942 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1888 LAYER M4 ;
  END BIAS_DBP[11]
  PIN BIAS_DBP[10] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.194 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.1856 LAYER M2 ;
  END BIAS_DBP[10]
  PIN BIAS_DBP[9] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.606 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9104 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.218 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.0032 LAYER M6 ;
  END BIAS_DBP[9]
  PIN BIAS_DBP[8] 
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
  END BIAS_DBP[8]
  PIN BIAS_DBP[7] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.029 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1716 LAYER M2 ;
  END BIAS_DBP[7]
  PIN BIAS_DBP[6] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
  END BIAS_DBP[6]
  PIN BIAS_DBP[5] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.982 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3648 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.966 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0944 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.398 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 50.1952 LAYER M6 ;
  END BIAS_DBP[5]
  PIN BIAS_DBP[4] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.692 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
  END BIAS_DBP[4]
  PIN BIAS_DBP[3] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.66 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.566 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.798 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1552 LAYER M4 ;
  END BIAS_DBP[3]
  PIN BIAS_DBP[2] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.618 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1632 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.898 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5952 LAYER M4 ;
  END BIAS_DBP[2]
  PIN BIAS_DBP[1] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.904 LAYER M3 ;
  END BIAS_DBP[1]
  PIN BIAS_DBP[0] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DBP[0]
  PIN BIAS_DBN[13] 
    ANTENNAPARTIALMETALAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.206 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M3 ;
  END BIAS_DBN[13]
  PIN BIAS_DBN[12] 
    ANTENNAPARTIALMETALAREA 0.0225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
  END BIAS_DBN[12]
  PIN BIAS_DBN[11] 
    ANTENNAPARTIALMETALAREA 0.031 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 3.124 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8336 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.218 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 18.6032 LAYER M6 ;
  END BIAS_DBN[11]
  PIN BIAS_DBN[10] 
    ANTENNAPARTIALMETALAREA 2.7495 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1418 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.426 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9184 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.958 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0592 LAYER M4 ;
  END BIAS_DBN[10]
  PIN BIAS_DBN[9] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.164 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1656 LAYER M3 ;
  END BIAS_DBN[9]
  PIN BIAS_DBN[8] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1562 LAYER M2 ;
  END BIAS_DBN[8]
  PIN BIAS_DBN[7] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
  END BIAS_DBN[7]
  PIN BIAS_DBN[6] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.802 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5728 LAYER M3 ;
  END BIAS_DBN[6]
  PIN BIAS_DBN[5] 
    ANTENNAPARTIALMETALAREA 0.048 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3608 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.482 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5648 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.062 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 44.3168 LAYER M6 ;
  END BIAS_DBN[5]
  PIN BIAS_DBN[4] 
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3608 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.104 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5016 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.678 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 38.2272 LAYER M6 ;
  END BIAS_DBN[4]
  PIN BIAS_DBN[3] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.702 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.578 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.618 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 29.1632 LAYER M6 ;
  END BIAS_DBN[3]
  PIN BIAS_DBN[2] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.338 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.0676 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.702 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.7328 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.878 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 30.3072 LAYER M6 ;
  END BIAS_DBN[2]
  PIN BIAS_DBN[1] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.724 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2736 LAYER M3 ;
  END BIAS_DBN[1]
  PIN BIAS_DBN[0] 
    ANTENNAPARTIALMETALAREA 0.4095 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8458 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.706 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1504 LAYER M3 ;
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13] 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.918 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0832 LAYER M3 ;
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9722 LAYER M2 ;
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10] 
    ANTENNAPARTIALMETALAREA 0.3885 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7534 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.618 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M3 ;
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.5805 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5982 LAYER M3 ;
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.822 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8608 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.838 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 43.3312 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 342.85 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1513.12 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0645 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3278 LAYER M2 ;
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.688 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.1152 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 5.638 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.8512 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.466 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 24.0944 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 97.0527 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 428.99 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA5 ;
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4] 
    ANTENNAPARTIALMETALAREA 0.358 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4384 LAYER M3 ;
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3] 
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0532 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.538 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 42.0112 LAYER M6 ;
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2] 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.242 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3088 LAYER M6 ;
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.446 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3608 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.578 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.7872 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.722 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 47.2208 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 291.853 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1287.19 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA6 ;
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.786 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.538 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0112 LAYER M4 ;
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13] 
    ANTENNAPARTIALMETALAREA 0.031 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M3 ;
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.165 LAYER M2 ;
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M4 ;
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.5825 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.007 LAYER M3 ;
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.456 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0504 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.266 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6144 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.158 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 31.5392 LAYER M6 ;
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.338 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.422 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9008 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.186 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2624 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.318 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 27.8432 LAYER M6 ;
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7552 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.458 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 28.4592 LAYER M6 ;
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.5195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.9298 LAYER M2 ;
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.158 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.3392 LAYER M4 ;
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1] 
    ANTENNAPARTIALMETALAREA 0.023 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1012 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.718 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6032 LAYER M3 ;
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0] 
    ANTENNAPARTIALMETALAREA 0.0195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.64 LAYER M3 ;
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.2455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0802 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M3 ;
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4] 
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.544 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8816 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.798 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5552 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 27.758 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 122.179 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 426.699 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1879.83 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA5 ;
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.091 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.5008 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 130.69 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.038 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.0112 LAYER M4 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 63.4675 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 280.877 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA4 ;
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.611 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7324 LAYER M2 ;
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.0665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.2524 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 182.505 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.1836 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 191.72 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.2165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9526 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.154 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1216 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.718 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 14.6573 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 65.8153 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA5 ;
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6112 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.791 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 82.7814 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.819672 LAYER VIA3 ;
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9458 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.786 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.6833 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 140.323 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.297 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.35 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.457 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.631 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.6128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.443 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 178.706 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.323625 LAYER VIA3 ;
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.632 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2248 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.9848 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 144.066 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[16] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.261 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1484 LAYER M2 ;
  END BIAS_TIA_G_POT[16]
  PIN BIAS_TIA_G_POT[15] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.198 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.5152 LAYER M3 ;
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14] 
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.6608 LAYER M3 ;
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13] 
    ANTENNAPARTIALMETALAREA 0.2255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9922 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.562 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 24.5168 LAYER M5 ;
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12] 
    ANTENNAPARTIALMETALAREA 0.181 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7964 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2992 LAYER M3 ;
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11] 
    ANTENNAPARTIALMETALAREA 1.0745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7278 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.942 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.3888 LAYER M3 ;
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1132 LAYER M2 ;
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.289 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3156 LAYER M2 ;
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.471 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0724 LAYER M2 ;
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7] 
    ANTENNAPARTIALMETALAREA 0.3325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M3 ;
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.994 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.406 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 60.518 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 266.323 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 12.538 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 55.2112 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 257.167 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1134.62 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5] 
    ANTENNAPARTIALMETALAREA 0.6255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7522 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.356 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.77092 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 44.7042 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4] 
    ANTENNAPARTIALMETALAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1132 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.19 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.68 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ; 
    ANTENNAMAXAREACAR 68.5417 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 304.825 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.0929 LAYER VIA4 ;
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.5425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.875 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.358 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.06818 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.5772 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.2886 LAYER VIA3 ;
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2] 
    ANTENNAPARTIALMETALAREA 0.187 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8228 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.382 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1248 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 49.5112 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 220.196 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA4 ;
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1] 
    ANTENNAPARTIALMETALAREA 0.3145 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3838 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M3 ;
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0] 
    ANTENNAPARTIALMETALAREA 0.051 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2244 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.946 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2064 LAYER M4 ;
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13] 
    ANTENNAPARTIALMETALAREA 0.123 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5412 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3 ;
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 7.988 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.3232 LAYER M2 ;
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.452 LAYER M2 ;
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.722 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0512 LAYER M4 ;
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6] 
    ANTENNAPARTIALMETALAREA 0.2245 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9878 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.4992 LAYER M4 ;
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5] 
    ANTENNAPARTIALMETALAREA 0.076 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.758 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3792 LAYER M3 ;
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.942 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1888 LAYER M3 ;
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3528 LAYER M2 ;
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2] 
    ANTENNAPARTIALMETALAREA 0.0195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M3 ;
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.039 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2156 LAYER M2 ;
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4158 LAYER M2 ;
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.8195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6058 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.7208 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 117.348 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.212 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3768 LAYER M2 ;
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7798 LAYER M2 ;
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.942 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1888 LAYER M4 ;
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.9225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.103 LAYER M2 ;
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.948 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1712 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.866 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.4913 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 84.961 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.5915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6026 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 71.7565 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 315.43 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA3 ;
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.537 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.626 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7984 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.718 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 74.7905 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 328.291 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA4 ;
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.4215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.6986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.618 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1632 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.4939 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.359 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA3 ;
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2] 
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.237 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0868 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.01 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.888 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 68.7925 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 304.155 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA4 ;
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.399 LAYER M2 ;
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.859 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7796 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.118 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9632 LAYER M3 ;
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.111 LAYER M2 ;
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.811 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.5178 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 183.896 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3 ;
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3298 LAYER M2 ;
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.138 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0512 LAYER M2 ;
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.4125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.747 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.806 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.918 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0832 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 65.4013 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 290.408 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA4 ;
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0] 
    ANTENNAPARTIALMETALAREA 1.153 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0732 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.87 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.6311 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 214.971 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.9885 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3934 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 LAYER M2 ; 
    ANTENNAMAXAREACAR 18.7589 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 82.3014 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.076 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8224 LAYER M3 ;
    ANTENNAGATEAREA 0.0564 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.8369 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 167.805 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.70922 LAYER VIA3 ;
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.586 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.184 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4976 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.106 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 20.662 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 90.9568 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 410.332 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1804.51 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA5 ;
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.126 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.938 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5712 LAYER M3 ;
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.55 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3232 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.532 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8288 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 19.278 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 84.8672 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1536 LAYER M5 ; 
    ANTENNAMAXAREACAR 140.603 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 618.307 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.520833 LAYER VIA5 ;
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.4755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0922 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3 ;
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.217 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9548 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.298 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M4 ;
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.998 LAYER M2 ;
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.8315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.6586 LAYER M2 ;
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0816 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.018 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5232 LAYER M4 ;
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.4985 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.2374 LAYER M2 ;
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.718 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M4 ;
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0512 LAYER M4 ;
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M3 ;
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1682 LAYER M2 ;
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.288 LAYER M2 ;
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4] 
    ANTENNAPARTIALMETALAREA 0.0705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3102 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7024 LAYER M3 ;
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.458 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0592 LAYER M4 ;
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3354 LAYER M2 ;
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1] 
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.802 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5728 LAYER M3 ;
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.165 LAYER M2 ;
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done 
    ANTENNAPARTIALMETALAREA 0.106 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4664 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.958 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.338 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.5312 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 1.678 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4272 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M7 ; 
    ANTENNAMAXAREACAR 193.875 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 853.402 LAYER M7 ;
    ANTENNAMAXCUTCAR 4.42804 LAYER VIA7 ;
  END dsadc_conv_done
  PIN dsadc_en 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.552 LAYER M2 ;
  END dsadc_en
  PIN dsadc_clk 
    ANTENNAPARTIALMETALAREA 1.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 65.384 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 72.0984 LAYER M3 ;
  END dsadc_clk
  PIN dsadc_switch[2] 
    ANTENNAPARTIALMETALAREA 0.347 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5268 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.5845 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0158 LAYER M3 ;
  END dsadc_switch[2]
  PIN dsadc_switch[1] 
    ANTENNAPARTIALMETALAREA 0.167 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7348 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.703 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1372 LAYER M3 ;
  END dsadc_switch[1]
  PIN dsadc_switch[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4762 LAYER M2 ;
  END dsadc_switch[0]
  PIN dac_en_pot 
    ANTENNAPARTIALMETALAREA 0.2245 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9878 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.646 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2864 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 4.142 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2688 LAYER M5 ;
  END dac_en_pot
  PIN adc_ext_in 
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.5568 LAYER M3 ;
  END adc_ext_in
  PIN atp_en 
    ANTENNAPARTIALMETALAREA 0.4445 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9558 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.8448 LAYER M3 ;
  END atp_en
  PIN atp_sel 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.357 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6148 LAYER M2 ;
  END atp_sel
  PIN adc_sel 
    ANTENNAPARTIALMETALAREA 0.0295 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.198 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.7152 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.206 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M4 ;
  END adc_sel
  PIN saradc_clk 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8534 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.4522 LAYER M3 ;
  END saradc_clk
  PIN saradc_rdy 
    ANTENNAPARTIALMETALAREA 0.3025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.331 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.378 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7072 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 11.078 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 48.7872 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M5 ; 
    ANTENNAMAXAREACAR 395.591 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1742.38 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.30548 LAYER VIA5 ;
  END saradc_rdy
  PIN saradc_rst 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.067 LAYER M2 ;
  END saradc_rst
  PIN saradc_data[9] 
    ANTENNAPARTIALMETALAREA 0.3115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3706 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 10.878 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 47.9072 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5 ; 
    ANTENNAMAXAREACAR 288.438 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1271.03 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.01511 LAYER VIA5 ;
  END saradc_data[9]
  PIN saradc_data[8] 
    ANTENNAPARTIALMETALAREA 0.4315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.338 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 58.7312 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 604.312 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2657.88 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[8]
  PIN saradc_data[7] 
    ANTENNAPARTIALMETALAREA 0.3555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6522 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M2 ; 
    ANTENNAMAXAREACAR 10.4484 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 46.9219 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.503778 LAYER VIA2 ;
  END saradc_data[7]
  PIN saradc_data[6] 
    ANTENNAPARTIALMETALAREA 0.187 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8228 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1815 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8426 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 9.898 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 43.5952 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.432 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6 ; 
    ANTENNAMAXAREACAR 58.5163 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 260.261 LAYER M6 ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6 ;
  END saradc_data[6]
  PIN saradc_data[5] 
    ANTENNAPARTIALMETALAREA 1.1625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.115 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.098 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8752 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.186 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 15.598 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 68.6752 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 689.537 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 3037.27 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[5]
  PIN saradc_data[4] 
    ANTENNAPARTIALMETALAREA 0.307 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.5615 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5146 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 12.858 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 56.6192 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 615.496 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2712.08 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[4]
  PIN saradc_data[3] 
    ANTENNAPARTIALMETALAREA 0.8425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.707 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.4048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 272.872 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1200.32 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END saradc_data[3]
  PIN saradc_data[2] 
    ANTENNAPARTIALMETALAREA 0.4425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2704 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 12.538 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 55.2112 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 586.027 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2580.36 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[2]
  PIN saradc_data[1] 
    ANTENNAPARTIALMETALAREA 0.5425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.387 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 14.738 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 64.8912 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 651.812 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2859.45 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.85714 LAYER VIA5 ;
  END saradc_data[1]
  PIN saradc_data[0] 
    ANTENNAPARTIALMETALAREA 0.9019 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7114 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.738 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6912 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.058 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.0992 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M6 ; 
    ANTENNAMAXAREACAR 183.685 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 813.94 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.267 LAYER VIA6 ;
  END saradc_data[0]
END MCU

END LIBRARY
