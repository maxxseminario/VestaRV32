

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO MCU 
  PIN resetn_in 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 25.782 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 113.485 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 974.013 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4292.32 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6 ;
  END resetn_in
  PIN resetn_out 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.474 LAYER M2 ;
  END resetn_out
  PIN resetn_dir 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6654 LAYER M2 ;
  END resetn_dir
  PIN resetn_ren 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1086 LAYER M2 ;
  END resetn_ren
  PIN prt1_in[7] 
    ANTENNAPARTIALMETALAREA 21.4525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 94.391 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.2928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 205.461 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 902.672 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt1_in[7]
  PIN prt1_in[6] 
    ANTENNAPARTIALMETALAREA 0.0805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0269 LAYER M2 ; 
    ANTENNAMAXAREACAR 91.0595 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 365.903 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.743494 LAYER VIA2 ;
  END prt1_in[6]
  PIN prt1_in[5] 
    ANTENNAPARTIALMETALAREA 1.5525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.831 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 7.108 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.3632 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 202.846 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 886.06 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END prt1_in[5]
  PIN prt1_in[4] 
    ANTENNAPARTIALMETALAREA 1.1525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.071 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.5968 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 514.887 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2265.91 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END prt1_in[4]
  PIN prt1_in[3] 
    ANTENNAPARTIALMETALAREA 0.176 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1936 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5862 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.976 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER M4 ; 
    ANTENNAMAXAREACAR 31.6541 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 42.2013 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.786164 LAYER VIA4 ;
  END prt1_in[3]
  PIN prt1_in[2] 
    ANTENNAPARTIALMETALAREA 2.1135 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3434 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.928 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.3712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 125.123 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 543.327 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[2]
  PIN prt1_in[1] 
    ANTENNAPARTIALMETALAREA 0.1755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7722 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.472 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.7648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 146.187 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 643.187 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[1]
  PIN prt1_in[0] 
    ANTENNAPARTIALMETALAREA 21.7355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 95.6362 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 LAYER M2 ; 
    ANTENNAMAXAREACAR 299.876 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 1317.2 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.271003 LAYER VIA2 ;
  END prt1_in[0]
  PIN prt1_out[7] 
    ANTENNAPARTIALMETALAREA 2.092 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2048 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.8528 LAYER M3 ;
  END prt1_out[7]
  PIN prt1_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.319 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.6916 LAYER M2 ;
  END prt1_out[6]
  PIN prt1_out[5] 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.4544 LAYER M3 ;
  END prt1_out[5]
  PIN prt1_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 8.121 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.7764 LAYER M2 ;
  END prt1_out[4]
  PIN prt1_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[3]
  PIN prt1_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.746 LAYER M2 ;
  END prt1_out[2]
  PIN prt1_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[1]
  PIN prt1_out[0] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
  END prt1_out[0]
  PIN prt1_dir[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[7]
  PIN prt1_dir[6] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
  END prt1_dir[6]
  PIN prt1_dir[5] 
    ANTENNAPARTIALMETALAREA 0.1165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3488 LAYER M3 ;
  END prt1_dir[5]
  PIN prt1_dir[4] 
    ANTENNAPARTIALMETALAREA 0.1965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8646 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.406 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M3 ;
  END prt1_dir[4]
  PIN prt1_dir[3] 
    ANTENNAPARTIALMETALAREA 1.4605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4262 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.0448 LAYER M3 ;
  END prt1_dir[3]
  PIN prt1_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.0425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.675 LAYER M2 ;
  END prt1_dir[2]
  PIN prt1_dir[1] 
    ANTENNAPARTIALMETALAREA 0.8915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9226 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
  END prt1_dir[1]
  PIN prt1_dir[0] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
  END prt1_dir[0]
  PIN prt1_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.4655 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.4922 LAYER M2 ;
  END prt1_ren[7]
  PIN prt1_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.3835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.9754 LAYER M2 ;
  END prt1_ren[6]
  PIN prt1_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.9635 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.9274 LAYER M2 ;
  END prt1_ren[5]
  PIN prt1_ren[4] 
    ANTENNAPARTIALMETALAREA 0.1075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.473 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.3008 LAYER M3 ;
  END prt1_ren[4]
  PIN prt1_ren[3] 
    ANTENNAPARTIALMETALAREA 0.2675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.177 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.086 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.2224 LAYER M3 ;
  END prt1_ren[3]
  PIN prt1_ren[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.3705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.3182 LAYER M2 ;
  END prt1_ren[2]
  PIN prt1_ren[1] 
    ANTENNAPARTIALMETALAREA 0.0475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.209 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
  END prt1_ren[1]
  PIN prt1_ren[0] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.209 LAYER M2 ;
  END prt1_ren[0]
  PIN prt2_in[7] 
    ANTENNAPARTIALMETALAREA 0.7735 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4474 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 LAYER M2 ; 
    ANTENNAMAXAREACAR 10.6222 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 45.187 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.185185 LAYER VIA2 ;
  END prt2_in[7]
  PIN prt2_in[6] 
    ANTENNAPARTIALMETALAREA 0.2975 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.353 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 13.0403 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 55.9539 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END prt2_in[6]
  PIN prt2_in[5] 
    ANTENNAPARTIALMETALAREA 0.7125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.135 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.55818 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 27.9858 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2 ;
  END prt2_in[5]
  PIN prt2_in[4] 
    ANTENNAPARTIALMETALAREA 0.7805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4782 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.58884 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 28.7594 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0786164 LAYER VIA2 ;
  END prt2_in[4]
  PIN prt2_in[3] 
    ANTENNAPARTIALMETALAREA 1.234 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5334 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.88784 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 9.43291 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.104822 LAYER VIA2 ;
  END prt2_in[3]
  PIN prt2_in[2] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 31.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 138.917 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 945.389 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4152.29 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt2_in[2]
  PIN prt2_in[1] 
    ANTENNAPARTIALMETALAREA 0.4555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0042 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 4.53774 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 19.0959 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2 ;
  END prt2_in[1]
  PIN prt2_in[0] 
    ANTENNAPARTIALMETALAREA 0.5305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3782 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.84067 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 16.3795 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.104822 LAYER VIA2 ;
  END prt2_in[0]
  PIN prt2_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.701 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1284 LAYER M2 ;
  END prt2_out[7]
  PIN prt2_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.681 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2 ;
  END prt2_out[6]
  PIN prt2_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.586 LAYER M2 ;
  END prt2_out[5]
  PIN prt2_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.737 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2868 LAYER M2 ;
  END prt2_out[4]
  PIN prt2_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.717 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1988 LAYER M2 ;
  END prt2_out[3]
  PIN prt2_out[2] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.514 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3056 LAYER M2 ;
  END prt2_out[2]
  PIN prt2_out[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.279 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2276 LAYER M2 ;
  END prt2_out[1]
  PIN prt2_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2 ;
  END prt2_out[0]
  PIN prt2_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7015 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1306 LAYER M2 ;
  END prt2_dir[7]
  PIN prt2_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1482 LAYER M2 ;
  END prt2_dir[6]
  PIN prt2_dir[5] 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.778 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.6672 LAYER M3 ;
  END prt2_dir[5]
  PIN prt2_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3486 LAYER M2 ;
  END prt2_dir[4]
  PIN prt2_dir[3] 
    ANTENNAPARTIALMETALAREA 0.731 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.9088 LAYER M3 ;
  END prt2_dir[3]
  PIN prt2_dir[2] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0218 LAYER M2 ;
  END prt2_dir[2]
  PIN prt2_dir[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0074 LAYER M2 ;
  END prt2_dir[1]
  PIN prt2_dir[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2254 LAYER M2 ;
  END prt2_dir[0]
  PIN prt2_ren[7] 
    ANTENNAPARTIALMETALAREA 0.6435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8314 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3808 LAYER M3 ;
  END prt2_ren[7]
  PIN prt2_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3166 LAYER M2 ;
  END prt2_ren[6]
  PIN prt2_ren[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.639 LAYER M2 ;
  END prt2_ren[5]
  PIN prt2_ren[4] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.409 LAYER M2 ;
  END prt2_ren[4]
  PIN prt2_ren[3] 
    ANTENNAPARTIALMETALAREA 0.6875 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.025 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.0368 LAYER M3 ;
  END prt2_ren[3]
  PIN prt2_ren[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5095 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2858 LAYER M2 ;
  END prt2_ren[2]
  PIN prt2_ren[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3095 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4058 LAYER M2 ;
  END prt2_ren[1]
  PIN prt2_ren[0] 
    ANTENNAPARTIALMETALAREA 0.4675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.057 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.2768 LAYER M3 ;
  END prt2_ren[0]
  PIN prt3_in[7] 
    ANTENNAPARTIALMETALAREA 24.0925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 106.007 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.6992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 419.631 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1846.08 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[7]
  PIN prt3_in[6] 
    ANTENNAPARTIALMETALAREA 16.2905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 71.7222 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 602.74 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2652.22 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2 ;
  END prt3_in[6]
  PIN prt3_in[5] 
    ANTENNAPARTIALMETALAREA 0.1725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.759 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.668 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.4272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 183.357 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 807.001 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.734684 LAYER VIA3 ;
  END prt3_in[5]
  PIN prt3_in[4] 
    ANTENNAPARTIALMETALAREA 0.6325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.783 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.814 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 52.1136 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 122.694 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 540.855 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
  END prt3_in[4]
  PIN prt3_in[3] 
    ANTENNAPARTIALMETALAREA 0.2355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0362 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.418 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.9712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 275.473 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1214.09 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 1.54769 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.338 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3312 LAYER M4 ;
    ANTENNAGATEAREA 0.1707 LAYER M4 ; 
    ANTENNAMAXAREACAR 289.17 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1274.61 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.54769 LAYER VIA4 ;
  END prt3_in[3]
  PIN prt3_in[2] 
    ANTENNAPARTIALMETALAREA 0.5755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4112 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M4 ; 
    ANTENNAMAXAREACAR 469.461 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 2052.69 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.21402 LAYER VIA4 ;
  END prt3_in[2]
  PIN prt3_in[1] 
    ANTENNAPARTIALMETALAREA 23.9155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 105.228 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.8288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 125.071 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 547.539 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.27669 LAYER VIA3 ;
  END prt3_in[1]
  PIN prt3_in[0] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 7.464 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.9296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 226.323 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 985.954 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt3_in[0]
  PIN prt3_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.803 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.2212 LAYER M2 ;
  END prt3_out[7]
  PIN prt3_out[6] 
    ANTENNAPARTIALMETALAREA 2.132 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4688 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.064 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.5696 LAYER M3 ;
  END prt3_out[6]
  PIN prt3_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.241 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1044 LAYER M2 ;
  END prt3_out[5]
  PIN prt3_out[4] 
    ANTENNAPARTIALMETALAREA 0.916 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0304 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.0608 LAYER M3 ;
  END prt3_out[4]
  PIN prt3_out[3] 
    ANTENNAPARTIALMETALAREA 3.612 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8928 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.046 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.8464 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.038 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6112 LAYER M4 ;
  END prt3_out[3]
  PIN prt3_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.996 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6704 LAYER M2 ;
  END prt3_out[2]
  PIN prt3_out[1] 
    ANTENNAPARTIALMETALAREA 1.392 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1248 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.928 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1712 LAYER M3 ;
  END prt3_out[1]
  PIN prt3_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.901 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2084 LAYER M2 ;
  END prt3_out[0]
  PIN prt3_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.2055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 62.5482 LAYER M2 ;
  END prt3_dir[7]
  PIN prt3_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.9615 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.9626 LAYER M2 ;
  END prt3_dir[6]
  PIN prt3_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt3_dir[5]
  PIN prt3_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
  END prt3_dir[4]
  PIN prt3_dir[3] 
    ANTENNAPARTIALMETALAREA 1.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6266 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.948 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.8592 LAYER M3 ;
  END prt3_dir[3]
  PIN prt3_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.3105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.5422 LAYER M2 ;
  END prt3_dir[2]
  PIN prt3_dir[1] 
    ANTENNAPARTIALMETALAREA 0.6515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.186 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M3 ;
  END prt3_dir[1]
  PIN prt3_dir[0] 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3 ;
  END prt3_dir[0]
  PIN prt3_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.3255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.7642 LAYER M2 ;
  END prt3_ren[7]
  PIN prt3_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.1235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6314 LAYER M2 ;
  END prt3_ren[6]
  PIN prt3_ren[5] 
    ANTENNAPARTIALMETALAREA 1.8385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1334 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.882 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5248 LAYER M3 ;
  END prt3_ren[5]
  PIN prt3_ren[4] 
    ANTENNAPARTIALMETALAREA 0.4405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9382 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.9888 LAYER M3 ;
  END prt3_ren[4]
  PIN prt3_ren[3] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.508 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.7232 LAYER M3 ;
  END prt3_ren[3]
  PIN prt3_ren[2] 
    ANTENNAPARTIALMETALAREA 11.8295 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 52.0938 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.8448 LAYER M3 ;
  END prt3_ren[2]
  PIN prt3_ren[1] 
    ANTENNAPARTIALMETALAREA 0.3675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4784 LAYER M3 ;
  END prt3_ren[1]
  PIN prt3_ren[0] 
    ANTENNAPARTIALMETALAREA 0.5405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M4 ;
  END prt3_ren[0]
  PIN prt4_in[7] 
    ANTENNAPARTIALMETALAREA 1.3555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9642 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 25.492 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 112.253 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 393.031 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1721.3 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.16802 LAYER VIA3 ;
  END prt4_in[7]
  PIN prt4_in[6] 
    ANTENNAPARTIALMETALAREA 2.4355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7162 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 18.638 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 82.1392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 301.336 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1328.07 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
  END prt4_in[6]
  PIN prt4_in[5] 
    ANTENNAPARTIALMETALAREA 1.2585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5374 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.246 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.7264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1456 LAYER M3 ; 
    ANTENNAMAXAREACAR 101.323 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 445.566 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.679368 LAYER VIA3 ;
  END prt4_in[5]
  PIN prt4_in[4] 
    ANTENNAPARTIALMETALAREA 4.1735 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.266 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 3.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2032 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 57.7228 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 256.328 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA4 ;
  END prt4_in[4]
  PIN prt4_in[3] 
    ANTENNAPARTIALMETALAREA 5.9505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.2262 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.3537 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.5488 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.734684 LAYER VIA3 ;
  END prt4_in[3]
  PIN prt4_in[2] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.284 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.1376 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1204 LAYER M3 ; 
    ANTENNAMAXAREACAR 244.321 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1073.69 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.16802 LAYER VIA3 ;
  END prt4_in[2]
  PIN prt4_in[1] 
    ANTENNAPARTIALMETALAREA 7.7685 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.2694 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M2 ; 
    ANTENNAMAXAREACAR 81.5253 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 356.295 LAYER M2 ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA2 ;
  END prt4_in[1]
  PIN prt4_in[0] 
    ANTENNAPARTIALMETALAREA 0.2725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 27.886 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 122.742 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 1080.52 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4736.44 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt4_in[0]
  PIN prt4_out[7] 
    ANTENNAPARTIALMETALAREA 8.492 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4006 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 70.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 77.264 LAYER M3 ;
  END prt4_out[7]
  PIN prt4_out[6] 
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 24.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.1062 LAYER M3 ;
  END prt4_out[6]
  PIN prt4_out[5] 
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.8502 LAYER M3 ;
  END prt4_out[5]
  PIN prt4_out[4] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0262 LAYER M3 ;
  END prt4_out[4]
  PIN prt4_out[3] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.1248 LAYER M3 ;
  END prt4_out[3]
  PIN prt4_out[2] 
    ANTENNAPARTIALMETALAREA 0.499 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1956 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.9024 LAYER M3 ;
  END prt4_out[2]
  PIN prt4_out[1] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.922 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 74.5008 LAYER M6 ;
  END prt4_out[1]
  PIN prt4_out[0] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[0]
  PIN prt4_dir[7] 
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.046 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.0464 LAYER M3 ;
  END prt4_dir[7]
  PIN prt4_dir[6] 
    ANTENNAPARTIALMETALAREA 0.651 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8644 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 15.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.4048 LAYER M3 ;
  END prt4_dir[6]
  PIN prt4_dir[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3222 LAYER M2 ;
  END prt4_dir[5]
  PIN prt4_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.2395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4538 LAYER M2 ;
  END prt4_dir[4]
  PIN prt4_dir[3] 
    ANTENNAPARTIALMETALAREA 0.871 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.118 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.5632 LAYER M3 ;
  END prt4_dir[3]
  PIN prt4_dir[2] 
    ANTENNAPARTIALMETALAREA 0.3565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5686 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.1328 LAYER M3 ;
  END prt4_dir[2]
  PIN prt4_dir[1] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 17.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 75.3808 LAYER M6 ;
  END prt4_dir[1]
  PIN prt4_dir[0] 
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6 ;
  END prt4_dir[0]
  PIN prt4_ren[7] 
    ANTENNAPARTIALMETALAREA 0.5475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.409 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.2448 LAYER M3 ;
  END prt4_ren[7]
  PIN prt4_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.497 LAYER M2 ;
  END prt4_ren[6]
  PIN prt4_ren[5] 
    ANTENNAPARTIALMETALAREA 1.1105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8862 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.266 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.2144 LAYER M3 ;
  END prt4_ren[5]
  PIN prt4_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.447 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3668 LAYER M2 ;
  END prt4_ren[4]
  PIN prt4_ren[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.2985 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7574 LAYER M2 ;
  END prt4_ren[3]
  PIN prt4_ren[2] 
    ANTENNAPARTIALMETALAREA 0.6835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.0448 LAYER M3 ;
  END prt4_ren[2]
  PIN prt4_ren[1] 
    ANTENNAPARTIALMETALAREA 0.8035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.342 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 71.9488 LAYER M6 ;
  END prt4_ren[1]
  PIN prt4_ren[0] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 17.146 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 75.4864 LAYER M6 ;
  END prt4_ren[0]
  PIN use_dac_glb_bias 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.3905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1182 LAYER M2 ;
  END use_dac_glb_bias
  PIN en_bias_buf 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1408 LAYER M2 ;
  END en_bias_buf
  PIN en_bias_gen 
    ANTENNAPARTIALMETALAREA 0.081 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.266 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M3 ;
  END en_bias_gen
  PIN BIAS_ADJ[5] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.566 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9344 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.918 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.8832 LAYER M6 ;
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.3465 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5686 LAYER M3 ;
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.067 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3388 LAYER M2 ;
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.856 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8544 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1664 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.178 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 44.8272 LAYER M6 ;
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
  END BIAS_DBP[13]
  PIN BIAS_DBP[12] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0655 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3322 LAYER M2 ;
  END BIAS_DBP[12]
  PIN BIAS_DBP[11] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.022 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.7408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.458 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.442 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3888 LAYER M5 ;
  END BIAS_DBP[11]
  PIN BIAS_DBP[10] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.6015 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0906 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.042 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6288 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 11.524 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 50.7936 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.968 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.684 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0976 LAYER M6 ;
  END BIAS_DBP[10]
  PIN BIAS_DBP[9] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.886 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5424 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.338 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.5312 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 331.127 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1460.58 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA6 ;
  END BIAS_DBP[9]
  PIN BIAS_DBP[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.2365 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4846 LAYER M2 ;
  END BIAS_DBP[8]
  PIN BIAS_DBP[7] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.778 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4672 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.358 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 32.4192 LAYER M6 ;
  END BIAS_DBP[7]
  PIN BIAS_DBP[6] 
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9152 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.426 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3184 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.498 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 37.4352 LAYER M6 ;
  END BIAS_DBP[6]
  PIN BIAS_DBP[5] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 7.776 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 34.3024 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.242 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9088 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 41.6108 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 186.069 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA5 ;
  END BIAS_DBP[5]
  PIN BIAS_DBP[4] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.398 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7952 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.906 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.8304 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.718 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 38.4032 LAYER M6 ;
  END BIAS_DBP[4]
  PIN BIAS_DBP[3] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.602 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6928 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.142 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8688 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.258 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 31.9792 LAYER M6 ;
  END BIAS_DBP[3]
  PIN BIAS_DBP[2] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.722 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.358 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.362 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0368 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.724 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.0736 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M6 ; 
    ANTENNAMAXAREACAR 166.391 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 737.28 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.23457 LAYER VIA6 ;
  END BIAS_DBP[2]
  PIN BIAS_DBP[1] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.882 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 39.1248 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 250.346 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1105.37 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA6 ;
  END BIAS_DBP[1]
  PIN BIAS_DBP[0] 
    ANTENNAPARTIALMETALAREA 0.0225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9152 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.606 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1104 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.894 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 52.4656 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 319.246 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1409.95 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6 ;
  END BIAS_DBP[0]
  PIN BIAS_DBN[13] 
    ANTENNAPARTIALMETALAREA 1.828 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0432 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6752 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.646 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2864 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.018 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.7232 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ; 
    ANTENNAMAXAREACAR 142.944 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 633.863 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.45902 LAYER VIA6 ;
  END BIAS_DBN[13]
  PIN BIAS_DBN[12] 
    ANTENNAPARTIALMETALAREA 0.0225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 5.016 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1584 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 2.238 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 9.8912 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 81.6414 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 360.799 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA6 ;
  END BIAS_DBN[12]
  PIN BIAS_DBN[11] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.644 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3216 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.018 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9232 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.258 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3792 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 91.3961 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 404.736 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_DBN[11]
  PIN BIAS_DBN[10] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9168 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.398 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1952 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.702 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.9328 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.74 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 29.744 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 157.627 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 697.165 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6 ;
  END BIAS_DBN[10]
  PIN BIAS_DBN[9] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.249 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0956 LAYER M2 ;
  END BIAS_DBN[9]
  PIN BIAS_DBN[8] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.338 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9312 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.946 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0064 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.338 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9312 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 140.256 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 619.085 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA6 ;
  END BIAS_DBN[8]
  PIN BIAS_DBN[7] 
    ANTENNAPARTIALMETALAREA 1.957 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6548 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.478 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.9472 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 153.82 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 679.799 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA4 ;
  END BIAS_DBN[7]
  PIN BIAS_DBN[6] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 179.269 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 789.443 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA3 ;
  END BIAS_DBN[6]
  PIN BIAS_DBN[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.698 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1152 LAYER M3 ;
  END BIAS_DBN[5]
  PIN BIAS_DBN[4] 
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.8848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.802 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1728 LAYER M6 ;
  END BIAS_DBN[4]
  PIN BIAS_DBN[3] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.738 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6912 LAYER M3 ;
  END BIAS_DBN[3]
  PIN BIAS_DBN[2] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.424 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M3 ; 
    ANTENNAMAXAREACAR 54.5813 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 233.704 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.823045 LAYER VIA3 ;
  END BIAS_DBN[2]
  PIN BIAS_DBN[1] 
    ANTENNAPARTIALMETALAREA 0.026 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1144 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.898 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9952 LAYER M4 ;
  END BIAS_DBN[1]
  PIN BIAS_DBN[0] 
    ANTENNAPARTIALMETALAREA 0.5165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2726 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M3 ;
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13] 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.078 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.5872 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.018 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9232 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.546 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2464 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.818 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.5312 LAYER M6 ;
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0245 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1518 LAYER M2 ;
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.328 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4032 LAYER M4 ;
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.498 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6352 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.198 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3152 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.178 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4272 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.968 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.498 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 41.8352 LAYER M6 ;
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.065 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.33 LAYER M2 ;
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8] 
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.538 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2112 LAYER M3 ;
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7] 
    ANTENNAPARTIALMETALAREA 0.119 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5676 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 30.712 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 123.183 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 544.39 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.666667 LAYER VIA4 ;
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.46 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.312 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 63.45 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 281.563 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA4 ;
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.731 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.9484 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.042 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.602 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4928 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 44.5274 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 196.609 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA4 ;
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4] 
    ANTENNAPARTIALMETALAREA 0.4275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.881 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.606 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1104 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.518 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.9232 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ; 
    ANTENNAMAXAREACAR 143.637 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 636.448 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.0929 LAYER VIA4 ;
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3] 
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.422 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.346 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9664 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.3 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.408 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 578.286 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2548.17 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.23625 LAYER VIA6 ;
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2] 
    ANTENNAPARTIALMETALAREA 0.7195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2098 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.66 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.402 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.104 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5016 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.238 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4912 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M6 ; 
    ANTENNAMAXAREACAR 103.493 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 458.16 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.85185 LAYER VIA6 ;
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1] 
    ANTENNAPARTIALMETALAREA 0.091 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.682 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 25.0448 LAYER M6 ;
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0] 
    ANTENNAPARTIALMETALAREA 0.0225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.398 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1952 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.548 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 37.7432 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 1.026 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5584 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 221.303 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 977.129 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA7 ;
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13] 
    ANTENNAPARTIALMETALAREA 0.457 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0548 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5808 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.018 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 30.9232 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ; 
    ANTENNAMAXAREACAR 259.539 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1147.62 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.18579 LAYER VIA6 ;
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.6675 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.381 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 3.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8512 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.968 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.358 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8192 LAYER M6 ;
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.338 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 32.3312 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 142.902 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 632.387 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA6 ;
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.122 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.7808 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.596 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 37.9104 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 181.058 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 800.498 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA6 ;
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.358 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8192 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.498 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.6352 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.968 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.622 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1808 LAYER M5 ;
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0928 LAYER M3 ;
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.582 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.578 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.7872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.146 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.978 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.7472 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 114.592 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 509.696 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.589 LAYER VIA6 ;
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.369 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6676 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.178 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2272 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.126 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M5 ; 
    ANTENNAMAXAREACAR 51.052 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 228.881 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.44033 LAYER VIA5 ;
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4] 
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.74 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.944 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ; 
    ANTENNAMAXAREACAR 142.914 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 621.454 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.63934 LAYER VIA4 ;
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.718 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.482 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.1648 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.782 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M5 ; 
    ANTENNAMAXAREACAR 25.0849 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 113.72 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.23457 LAYER VIA5 ;
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.398 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7952 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.318 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.6432 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.326 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4784 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M5 ; 
    ANTENNAMAXAREACAR 64.2207 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 285.918 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.23457 LAYER VIA5 ;
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6148 LAYER M3 ;
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.9655 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2482 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.942 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1888 LAYER M3 ;
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.556 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.142 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0688 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 28.958 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 127.459 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.182 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4448 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 97.1537 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 426.814 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3] 
    ANTENNAPARTIALMETALAREA 1.1175 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.917 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M3 ;
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.232 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.402 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2128 LAYER M4 ;
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.278 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M2 ;
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.35 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.54 LAYER M2 ;
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.2555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M3 ;
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.269 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6276 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.518 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7232 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ; 
    ANTENNAMAXAREACAR 76.6189 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 337.978 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.63934 LAYER VIA4 ;
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.1845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8118 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.042 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.878 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9072 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.354 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0016 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 23.373 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 104.165 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA5 ;
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.271 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.648 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3392 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 34.1378 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 151.887 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA5 ;
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.2975 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.309 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.368 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.0546 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 177.709 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0] 
    ANTENNAPARTIALMETALAREA 0.043 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.308 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8432 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 70.3644 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 311.96 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.7316 LAYER VIA5 ;
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[15] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.9775 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.301 LAYER M2 ;
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14] 
    ANTENNAPARTIALMETALAREA 0.123 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5412 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.438 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9712 LAYER M3 ;
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13] 
    ANTENNAPARTIALMETALAREA 0.027 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1188 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.962 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 26.2768 LAYER M5 ;
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12] 
    ANTENNAPARTIALMETALAREA 0.157 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6908 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.702 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1328 LAYER M4 ;
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3386 LAYER M2 ;
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10] 
    ANTENNAPARTIALMETALAREA 0.187 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8228 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.288 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3112 LAYER M3 ;
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9] 
    ANTENNAPARTIALMETALAREA 0.3635 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5994 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.418 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M3 ;
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.288 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3 ;
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1318 LAYER M2 ;
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.709 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1636 LAYER M2 ;
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5] 
    ANTENNAPARTIALMETALAREA 0.6255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7522 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.436 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.2529 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.6248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.626 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7984 LAYER M4 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 21.2861 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 96.0058 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.438 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9712 LAYER M5 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 27.6064 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 124.45 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA5 ;
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4] 
    ANTENNAPARTIALMETALAREA 1.471 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4724 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.2821 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 170.481 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.819672 LAYER VIA3 ;
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3295 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4938 LAYER M2 ;
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2] 
    ANTENNAPARTIALMETALAREA 0.353 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5532 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.206 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M4 ;
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9742 LAYER M2 ;
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.713 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1812 LAYER M2 ;
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13] 
    ANTENNAPARTIALMETALAREA 0.282 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.898 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7952 LAYER M4 ;
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3 ;
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.458 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0592 LAYER M3 ;
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.998 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4352 LAYER M4 ;
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.318 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4432 LAYER M3 ;
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.026 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1584 LAYER M2 ;
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7766 LAYER M2 ;
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.142 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M3 ;
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6928 LAYER M3 ;
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.846 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7664 LAYER M3 ;
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2] 
    ANTENNAPARTIALMETALAREA 0.0825 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.363 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.626 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7984 LAYER M3 ;
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.179 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8316 LAYER M2 ;
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0] 
    ANTENNAPARTIALMETALAREA 0.0395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1738 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3 ;
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.111 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4884 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0635 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3234 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.31 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.208 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 36.0426 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 159.276 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4 ;
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.214 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9416 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.778 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4672 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.802 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 27.702 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 121.933 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 3.346 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7664 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M7 ; 
    ANTENNAMAXAREACAR 149.549 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 660.332 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.7316 LAYER VIA7 ;
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.1245 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5478 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.102 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8928 LAYER M4 ;
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.758 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3352 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 12.2042 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 52.2049 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.9545 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 56.1414 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.906 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0304 LAYER M4 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 26.0281 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 114.3 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA4 ;
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.431 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8964 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9568 LAYER M3 ;
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.271 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.071 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3564 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.962 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6768 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 45.956 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 203.518 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA4 ;
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.7915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4826 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1008 LAYER M3 ;
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.034 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.6128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 100.357 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 441.482 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA3 ;
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.5265 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3166 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.336 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.7468 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 223.431 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.247 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0868 LAYER M2 ;
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.111 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4884 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.338 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.302 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7728 LAYER M4 ;
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 1.063 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6772 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.222 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.598 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 29.0752 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 3.582 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8048 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 LAYER M7 ; 
    ANTENNAMAXAREACAR 97.9587 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 431.279 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA7 ;
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.9685 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2614 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.686 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0624 LAYER M3 ;
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4] 
    ANTENNAPARTIALMETALAREA 1.385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.138 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.218 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.8032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.166 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 51.9385 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 231.172 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA4 ;
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.3805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6742 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.7328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.33 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.296 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 39.9657 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 177.561 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4 ;
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.133 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5852 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.036 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.4464 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 113.621 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 504 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA4 ;
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.0665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.586 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M5 ; 
    ANTENNAMAXAREACAR 182.1 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 805.307 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.26537 LAYER VIA5 ;
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.645 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.282 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.30097 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 28.7184 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.7785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4254 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.986 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3824 LAYER M3 ;
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4] 
    ANTENNAPARTIALMETALAREA 1.517 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6748 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.984 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.226 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 21.498 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 94.6352 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 1.906 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4304 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 124.093 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 542.061 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA7 ;
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3] 
    ANTENNAPARTIALMETALAREA 1.1505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0622 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.902 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M3 ; 
    ANTENNAMAXAREACAR 63.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 280.305 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.823045 LAYER VIA3 ;
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.587 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5828 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.708 LAYER M3 ;
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.351 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5088 LAYER M3 ;
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.674 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9656 LAYER M2 ;
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13] 
    ANTENNAPARTIALMETALAREA 4.553 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.1212 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.858 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8192 LAYER M4 ;
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.7135 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.1834 LAYER M2 ;
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.086 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.4224 LAYER M2 ;
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0816 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.536 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2464 LAYER M4 ;
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9] 
    ANTENNAPARTIALMETALAREA 1.295 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.646 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8864 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.658 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3392 LAYER M4 ;
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8] 
    ANTENNAPARTIALMETALAREA 0.0695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3058 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9632 LAYER M4 ;
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6] 
    ANTENNAPARTIALMETALAREA 0.1385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6094 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.378 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7072 LAYER M4 ;
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0855 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4202 LAYER M2 ;
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.642 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8688 LAYER M3 ;
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2] 
    ANTENNAPARTIALMETALAREA 0.0765 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3366 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.022 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5408 LAYER M3 ;
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1] 
    ANTENNAPARTIALMETALAREA 0.071 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3124 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.062 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7168 LAYER M3 ;
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0] 
    ANTENNAPARTIALMETALAREA 0.586 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.646 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8864 LAYER M3 ;
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done 
    ANTENNAPARTIALMETALAREA 0.625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.75 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.2608 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M3 ; 
    ANTENNAMAXAREACAR 519.306 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2286.91 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.22449 LAYER VIA3 ;
  END dsadc_conv_done
  PIN dsadc_en 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.141 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6644 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.398 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7952 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.062 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.3168 LAYER M5 ;
  END dsadc_en
  PIN dsadc_clk 
    ANTENNAPARTIALMETALAREA 0.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0934 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.624 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7624 LAYER M3 ;
  END dsadc_clk
  PIN dsadc_switch[2] 
    ANTENNAPARTIALMETALAREA 0.0895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3938 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1808 LAYER M3 ;
  END dsadc_switch[2]
  PIN dsadc_switch[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.358 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M2 ;
  END dsadc_switch[1]
  PIN dsadc_switch[0] 
    ANTENNAPARTIALMETALAREA 0.4385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9294 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.546 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4464 LAYER M3 ;
  END dsadc_switch[0]
  PIN dac_en_pot 
    ANTENNAPARTIALMETALAREA 0.0665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.086 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4224 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.858 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0192 LAYER M5 ;
  END dac_en_pot
  PIN adc_ext_in 
    ANTENNAPARTIALMETALAREA 0.451 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9844 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.698 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.1152 LAYER M3 ;
  END adc_ext_in
  PIN atp_en 
    ANTENNAPARTIALMETALAREA 0.3025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.375 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.738 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6912 LAYER M5 ;
  END atp_en
  PIN atp_sel 
    ANTENNAPARTIALMETALAREA 0.891 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9204 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.078 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.3872 LAYER M3 ;
  END atp_sel
  PIN adc_sel 
    ANTENNAPARTIALMETALAREA 0.6925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.047 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.0128 LAYER M3 ;
  END adc_sel
  PIN saradc_clk 
    ANTENNAPARTIALMETALAREA 3.162 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.642 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8822 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.576 LAYER M4 ;
  END saradc_clk
  PIN saradc_rdy 
    ANTENNAPARTIALMETALAREA 0.209 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9636 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.492 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.138 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 3.598 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8752 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M7 ; 
    ANTENNAMAXAREACAR 318.703 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 1407.83 LAYER M7 ;
    ANTENNAMAXCUTCAR 3.45821 LAYER VIA7 ;
  END saradc_rdy
  PIN saradc_rst 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1726 LAYER M2 ;
  END saradc_rst
  PIN saradc_data[9] 
    ANTENNAPARTIALMETALAREA 0.8865 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9006 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.638 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.4512 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.104 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5016 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 7.098 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 31.2752 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5 ; 
    ANTENNAMAXAREACAR 201.698 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 889.768 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.51134 LAYER VIA5 ;
  END saradc_data[9]
  PIN saradc_data[8] 
    ANTENNAPARTIALMETALAREA 0.2425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.067 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.546 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4464 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 17.918 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 78.8832 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M5 ; 
    ANTENNAMAXAREACAR 539.951 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2379.8 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.01729 LAYER VIA5 ;
  END saradc_data[8]
  PIN saradc_data[7] 
    ANTENNAPARTIALMETALAREA 0.7115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1306 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.766 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.2144 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 12.618 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 55.5632 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M5 ; 
    ANTENNAMAXAREACAR 411.037 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1809.7 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.30548 LAYER VIA5 ;
  END saradc_data[7]
  PIN saradc_data[6] 
    ANTENNAPARTIALMETALAREA 0.2665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1726 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.378 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5072 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.426 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9184 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.018 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5232 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.106 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 2.502 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 11.0528 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M7 ; 
    ANTENNAMAXAREACAR 438.772 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 1927.26 LAYER M7 ;
    ANTENNAMAXCUTCAR 3.45821 LAYER VIA7 ;
  END saradc_data[6]
  PIN saradc_data[5] 
    ANTENNAPARTIALMETALAREA 0.391 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7204 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.9395 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.2218 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 462.069 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2035.85 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.864553 LAYER VIA3 ;
  END saradc_data[5]
  PIN saradc_data[4] 
    ANTENNAPARTIALMETALAREA 0.4825 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.123 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 7.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.1552 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 7.516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 33.1584 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M5 ; 
    ANTENNAMAXAREACAR 230.346 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1017.38 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.30548 LAYER VIA5 ;
  END saradc_data[4]
  PIN saradc_data[3] 
    ANTENNAPARTIALMETALAREA 0.4915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1626 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.538 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.398 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 58.9952 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M5 ; 
    ANTENNAMAXAREACAR 417.965 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1833.38 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.30548 LAYER VIA5 ;
  END saradc_data[3]
  PIN saradc_data[2] 
    ANTENNAPARTIALMETALAREA 0.3055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.818 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.0836 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 185.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END saradc_data[2]
  PIN saradc_data[1] 
    ANTENNAPARTIALMETALAREA 0.8955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9402 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.1344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.458 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.2592 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.106 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 1.198 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3152 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M7 ; 
    ANTENNAMAXAREACAR 580.312 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 2554.11 LAYER M7 ;
    ANTENNAMAXCUTCAR 4.89796 LAYER VIA7 ;
  END saradc_data[1]
  PIN saradc_data[0] 
    ANTENNAPARTIALMETALAREA 0.8515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7466 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.438 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3712 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.106 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.338 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3312 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 2.082 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2048 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0269 LAYER M7 ; 
    ANTENNAMAXAREACAR 474.996 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 2081.39 LAYER M7 ;
    ANTENNAMAXCUTCAR 4.46097 LAYER VIA7 ;
  END saradc_data[0]
END MCU

END LIBRARY
