#******
# TECH LIB NAME: tsmc065
#
# The R,C and thickness values used in this LEF are typical values.
# These are taken from the
#   
# Document Title : TSMC 65NM CMOS LOGIC LOW POWER 1P9M SALICIDE CU_LOWK
#                  1.2 & 2.5V HD BEOL SPICE MODEL (CLN65LP)
# Document No    : T-N65-CL-SP-009 Version 1.1 03/09/2006.
#  
# DESIGN RULES ARE TAKEN FROM THE DOCUMENT
#
# Document Title : TSMC 65NM CMOS LOGIC DESIGN RULES
# Document No    : T-N65-CL-DR-001 Version 1.2 Apr 14, 2006. 
#
# Resistance and Capacitance Values
# ---------------------------------
# The LEF technology files included in this directory contain resistance and
# capacitance (RC) values for the purpose of timing driven place & route.
# Please note that the RC values contained in this tech file were created using
# the worst case interconnect models from the foundry and assume a full metal
# route at every grid location on every metal layer, so the values are
# intentionally very conservative. It is assumed that this technology file will
# be used only as a starting point for creating initial timing driven place &
# route runs during the development of your own more accurate RC values,
# tailored to your specific place & route environment. AS A RESULT, TIMING
# NUMBERS DERIVED FROM THESE RC VALUES MAY BE SIGNIFICANTLY SLOWER THAN
# REALITY.
# 
# The RC values used in the LEF technology file are to be used only for timing
# driven place & route. Due to accuracy limitations, please do not attempt to
# use this file for chip-level RC extraction in conjunction with your sign-off
# timing simulations. For chip-level extraction, please use a dedicated
# extraction tool such as HyperExtract, starRC or Fire & Ice QX, etc.
#
# Antenna Effect Properties
# -------------------------
# Antenna effect properties were modeled based on the following design rule
# document:
#
# Document No. T-N65-CL-DR-001 (TSMC 65NM CMOS LOGIC DESIGN RULE
#                            Version 1.2 04/14/2006 )
#
# $Id: tsmc_cln65_6X1Z_tech.lef,v 1.1 2006/12/26 09:02:36 pmullur Exp $
#
#******
VERSION 5.6 ;
# NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;

UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;
USEMINSPACING PIN OFF ;
USEMINSPACING OBS OFF ;

PROPERTYDEFINITIONS
    LAYER LEF57_SPACING STRING  ;
    LAYER LEF57_MINSTEP STRING ;
END PROPERTYDEFINITIONS

LAYER RVT
    TYPE IMPLANT ;
    WIDTH 0.18 ;
    SPACING 0.18 ;
END RVT

LAYER HVT
    TYPE IMPLANT ;
    WIDTH 0.18 ;
    SPACING 0.18 ;
END HVT 

LAYER LVT
    TYPE IMPLANT ;
    WIDTH 0.18 ;
    SPACING 0.18 ;
END LVT 

LAYER POLY1
    TYPE MASTERSLICE ;
END POLY1

LAYER M1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.20 ;
    OFFSET 0.10 ;
    WIDTH 0.09 ;
    MAXWIDTH 12.00 ; 
    AREA 0.042 ;
    SPACINGTABLE
    PARALLELRUNLENGTH 0.00 0.38 0.42 1.50 4.50
    WIDTH 0.00        0.09 0.09 0.09 0.09 0.09
    WIDTH 0.20        0.09 0.11 0.11 0.11 0.11
    WIDTH 0.42        0.09 0.11 0.16 0.16 0.16
    WIDTH 1.50        0.09 0.11 0.16 0.50 0.50
    WIDTH 4.50        0.09 0.11 0.16 0.50 1.50 ;
    MINENCLOSEDAREA  0.20 ;
    PROPERTY LEF57_MINSTEP "MINSTEP 0.09 MAXEDGES 1 ;" ;
    PROPERTY LEF57_SPACING "SPACING 0.11 ENDOFLINE 0.11 WITHIN 0.035 PARALLELEDGE 0.11 WITHIN 0.11 ;" ;
    MINIMUMCUT 2 WIDTH 0.30 ;
    MINIMUMCUT 4 WIDTH 0.70 ;
    MINIMUMCUT 2 WIDTH 0.3 LENGTH  0.3 WITHIN 0.8 ;
    MINIMUMCUT 2 WIDTH 2.0 LENGTH  2.0 WITHIN 2 ;
    MINIMUMCUT 2 WIDTH 3.0 LENGTH 10.0 WITHIN 5 ;
    ANTENNACUMAREARATIO 4996 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 4996 ) ( 0.059 4996 ) ( 0.06 43017 ) ( 1 43436 ) ) ;
    THICKNESS 0.18 ;
    HEIGHT 0.29 ;
    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
    FILLACTIVESPACING 0.61 ;
    RESISTANCE RPERSQ       1.6000e-01 ;
    CAPACITANCE CPERSQDIST  3.6364e-04 ;
    EDGECAPACITANCE        10.4194e-05 ;
END M1

LAYER VIA1
    TYPE CUT ;
    SPACING 0.13 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    ENCLOSURE BELOW 0.04 0.00 ;
    ENCLOSURE ABOVE 0.04 0.00 ;
    PREFERENCLOSURE BELOW 0.07 0.00 ;
    PREFERENCLOSURE ABOVE 0.07 0.00 ;
    ANTENNAAREARATIO 19 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 19 ) ( 0.059 19 ) ( 0.06 903 ) ( 1 1098 ) ) ;
END VIA1

LAYER M2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.20 ;
    OFFSET 0.10 ; 
    WIDTH 0.10 ;
    MAXWIDTH 12.00 ; 
    AREA 0.052 ;
    SPACINGTABLE
    PARALLELRUNLENGTH 0.00 0.38 0.40 1.50 4.50
    WIDTH 0.00        0.10 0.10 0.10 0.10 0.10
    WIDTH 0.20        0.10 0.12 0.12 0.12 0.12
    WIDTH 0.40        0.10 0.12 0.16 0.16 0.16
    WIDTH 1.50        0.10 0.12 0.16 0.50 0.50     
    WIDTH 4.50        0.10 0.12 0.16 0.50 1.50 ;
    MINENCLOSEDAREA  0.20 ;
    PROPERTY LEF57_MINSTEP "MINSTEP 0.10 MAXEDGES 1 ;" ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    MINIMUMCUT 2 WIDTH 0.30 ;
    MINIMUMCUT 4 WIDTH 0.70 ;
    MINIMUMCUT 2 WIDTH 0.3 LENGTH  0.3 WITHIN 0.8 ;
    MINIMUMCUT 2 WIDTH 2.0 LENGTH  2.0 WITHIN 2 ;
    MINIMUMCUT 2 WIDTH 3.0 LENGTH 10.0 WITHIN 5 ;
    ANTENNACUMAREARATIO 4996 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 4996 ) ( 0.059 4996 ) ( 0.06 43017 ) ( 1 43436 ) ) ;
    THICKNESS 0.22 ;
    HEIGHT 0.645 ;
    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
    FILLACTIVESPACING 0.61 ;
    RESISTANCE RPERSQ       1.4000e-01 ;
    CAPACITANCE CPERSQDIST  4.6607e-04 ;
    EDGECAPACITANCE        10.0799e-05 ;
END M2

LAYER VIA2
    TYPE CUT ;
    SPACING 0.13 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    ENCLOSURE BELOW 0.04 0.00 ;
    ENCLOSURE ABOVE 0.04 0.00 ;
    PREFERENCLOSURE BELOW 0.07 0.00 ;
    PREFERENCLOSURE ABOVE 0.07 0.00 ;
    ANTENNAAREARATIO 19 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 19 ) ( 0.059 19 ) ( 0.06 903 ) ( 1 1098 ) ) ;
END VIA2

LAYER M3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.20 ;
    OFFSET 0.10 ;
    WIDTH 0.10 ;
    MAXWIDTH 12.00 ; 
    AREA 0.052 ;
    SPACINGTABLE
    PARALLELRUNLENGTH 0.00 0.38 0.40 1.50 4.50
    WIDTH 0.00        0.10 0.10 0.10 0.10 0.10
    WIDTH 0.20        0.10 0.12 0.12 0.12 0.12
    WIDTH 0.40        0.10 0.12 0.16 0.16 0.16
    WIDTH 1.50        0.10 0.12 0.16 0.50 0.50     
    WIDTH 4.50        0.10 0.12 0.16 0.50 1.50 ;
    MINENCLOSEDAREA  0.20 ;
    PROPERTY LEF57_MINSTEP "MINSTEP 0.10 MAXEDGES 1 ;" ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    MINIMUMCUT 2 WIDTH 0.30 ;
    MINIMUMCUT 4 WIDTH 0.70 ;
    MINIMUMCUT 2 WIDTH 0.3 LENGTH  0.3 WITHIN 0.8 ;
    MINIMUMCUT 2 WIDTH 2.0 LENGTH  2.0 WITHIN 2 ;
    MINIMUMCUT 2 WIDTH 3.0 LENGTH 10.0 WITHIN 5 ;
    ANTENNACUMAREARATIO 4996 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 4996 ) ( 0.059 4996 ) ( 0.06 43017 ) ( 1 43436 ) ) ;
    THICKNESS 0.22 ;
    HEIGHT 1.04 ;
    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
    FILLACTIVESPACING 0.61 ;
    RESISTANCE RPERSQ       1.4000e-01 ;
    CAPACITANCE CPERSQDIST  4.6700e-04 ;
    EDGECAPACITANCE        10.1472e-05 ;
END M3

LAYER VIA3
    TYPE CUT ;
    SPACING 0.13 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    ENCLOSURE BELOW 0.04 0.00 ;
    ENCLOSURE ABOVE 0.04 0.00 ;
    PREFERENCLOSURE BELOW 0.07 0.00 ;
    PREFERENCLOSURE ABOVE 0.07 0.00 ;
    ANTENNAAREARATIO 19 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 19 ) ( 0.059 19 ) ( 0.06 903 ) ( 1 1098 ) ) ;
END VIA3

LAYER M4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    WIDTH 0.10 ;
    MAXWIDTH 12.00 ; 
    PITCH 0.20 ;
    OFFSET 0.10 ;
    AREA 0.052 ;
    SPACINGTABLE
    PARALLELRUNLENGTH 0.00 0.38 0.40 1.50 4.50
    WIDTH 0.00        0.10 0.10 0.10 0.10 0.10
    WIDTH 0.20        0.10 0.12 0.12 0.12 0.12
    WIDTH 0.40        0.10 0.12 0.16 0.16 0.16
    WIDTH 1.50        0.10 0.12 0.16 0.50 0.50     
    WIDTH 4.50        0.10 0.12 0.16 0.50 1.50 ;
    MINENCLOSEDAREA  0.20 ;
    PROPERTY LEF57_MINSTEP "MINSTEP 0.10 MAXEDGES 1 ;" ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    MINIMUMCUT 2 WIDTH 0.30 ;
    MINIMUMCUT 4 WIDTH 0.70 ;
    MINIMUMCUT 2 WIDTH 0.3 LENGTH  0.3 WITHIN 0.8 ;
    MINIMUMCUT 2 WIDTH 2.0 LENGTH  2.0 WITHIN 2 ;
    MINIMUMCUT 2 WIDTH 3.0 LENGTH 10.0 WITHIN 5 ;
    ANTENNACUMAREARATIO 4996 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 4996 ) ( 0.059 4996 ) ( 0.06 43017 ) ( 1 43436 ) ) ;
    THICKNESS 0.22 ;
    HEIGHT 1.435 ;
    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
    FILLACTIVESPACING 0.61 ;
    RESISTANCE RPERSQ       1.4000e-01 ;
    CAPACITANCE CPERSQDIST  4.6700e-04 ;
    EDGECAPACITANCE        10.1472e-05 ;
END M4

LAYER VIA4
    TYPE CUT ;
    SPACING 0.13 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    ENCLOSURE BELOW 0.04 0.00 ;
    ENCLOSURE ABOVE 0.04 0.00 ;
    PREFERENCLOSURE BELOW 0.07 0.00 ;
    PREFERENCLOSURE ABOVE 0.07 0.00 ;
    ANTENNAAREARATIO 19 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 19 ) ( 0.059 19 ) ( 0.06 903 ) ( 1 1098 ) ) ;
END VIA4

LAYER M5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.10 ;
    MAXWIDTH 12.00 ; 
    PITCH 0.20 ;
    OFFSET 0.10 ;
    AREA 0.052 ;
    SPACINGTABLE
    PARALLELRUNLENGTH 0.00 0.38 0.40 1.50 4.50
    WIDTH 0.00        0.10 0.10 0.10 0.10 0.10
    WIDTH 0.20        0.10 0.12 0.12 0.12 0.12
    WIDTH 0.40        0.10 0.12 0.16 0.16 0.16
    WIDTH 1.50        0.10 0.12 0.16 0.50 0.50     
    WIDTH 4.50        0.10 0.12 0.16 0.50 1.50 ;
    MINENCLOSEDAREA  0.20 ;
    PROPERTY LEF57_MINSTEP "MINSTEP 0.10 MAXEDGES 1 ;" ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    MINIMUMCUT 2 WIDTH 0.30 ;
    MINIMUMCUT 4 WIDTH 0.70 ;
    MINIMUMCUT 2 WIDTH 0.3 LENGTH  0.3 WITHIN 0.8 ;
    MINIMUMCUT 2 WIDTH 2.0 LENGTH  2.0 WITHIN 2 ;
    MINIMUMCUT 2 WIDTH 3.0 LENGTH 10.0 WITHIN 5 ;
    ANTENNACUMAREARATIO 4996 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 4996 ) ( 0.059 4996 ) ( 0.06 43017 ) ( 1 43436 ) ) ;
    THICKNESS 0.22 ;
    HEIGHT 1.83 ;
    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
    FILLACTIVESPACING 0.61 ;
    RESISTANCE RPERSQ      1.4000e-01 ;
    CAPACITANCE CPERSQDIST  4.6700e-04 ;
    EDGECAPACITANCE        10.1472e-05 ;
END M5

LAYER VIA5
    TYPE CUT ;
    SPACING 0.13 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    ENCLOSURE BELOW 0.04 0.00 ;
    ENCLOSURE ABOVE 0.04 0.00 ;
    PREFERENCLOSURE BELOW 0.07 0.00 ;
    PREFERENCLOSURE ABOVE 0.07 0.00 ;
    ANTENNAAREARATIO 19 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 19 ) ( 0.059 19 ) ( 0.06 903 ) ( 1 1098 ) ) ;
END VIA5

LAYER M6
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    WIDTH 0.10 ;
    MAXWIDTH 12.00 ; 
    PITCH 0.20 ;
    OFFSET 0.10 ;
    AREA 0.052 ;
    SPACINGTABLE
    PARALLELRUNLENGTH 0.00 0.38 0.40 1.50 4.50
    WIDTH 0.00        0.10 0.10 0.10 0.10 0.10
    WIDTH 0.20        0.10 0.12 0.12 0.12 0.12
    WIDTH 0.40        0.10 0.12 0.16 0.16 0.16
    WIDTH 1.50        0.10 0.12 0.16 0.50 0.50     
    WIDTH 4.50        0.10 0.12 0.16 0.50 1.50 ;
    MINENCLOSEDAREA  0.20 ;
    PROPERTY LEF57_MINSTEP "MINSTEP 0.10 MAXEDGES 1 ;" ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    MINIMUMCUT 2 WIDTH 0.30 ;
    MINIMUMCUT 4 WIDTH 0.70 ;
    MINIMUMCUT 2 WIDTH 0.3 LENGTH  0.3 WITHIN 0.8 ;
    MINIMUMCUT 2 WIDTH 2.0 LENGTH  2.0 WITHIN 2 ;
    MINIMUMCUT 2 WIDTH 3.0 LENGTH 10.0 WITHIN 5 ;
    ANTENNACUMAREARATIO 4996 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 4996 ) ( 0.059 4996 ) ( 0.06 43017 ) ( 1 43436 ) ) ;
    THICKNESS 0.22 ;
    HEIGHT 2.225 ;
    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
    FILLACTIVESPACING 0.61 ;
    RESISTANCE RPERSQ       1.4000e-01 ;
    CAPACITANCE CPERSQDIST  4.5882e-04 ;
    EDGECAPACITANCE        10.1038e-05 ;
END M6

LAYER VIA6
    TYPE CUT ;
    SPACING 0.13 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    ENCLOSURE BELOW 0.04 0.00 ;
    ENCLOSURE ABOVE 0.04 0.00 ;
    PREFERENCLOSURE BELOW 0.07 0.00 ;
    PREFERENCLOSURE ABOVE 0.07 0.00 ;
    ANTENNAAREARATIO 19 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 19 ) ( 0.059 19 ) ( 0.06 903 ) ( 1 1098 ) ) ;
END VIA6

LAYER M7
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.10 ;
    MAXWIDTH 12.00 ; 
    PITCH 0.20 ;
    OFFSET 0.10 ;
    AREA 0.052 ;
    SPACINGTABLE
    PARALLELRUNLENGTH 0.00 0.38 0.40 1.50 4.50
    WIDTH 0.00        0.10 0.10 0.10 0.10 0.10
    WIDTH 0.20        0.10 0.12 0.12 0.12 0.12
    WIDTH 0.40        0.10 0.12 0.16 0.16 0.16
    WIDTH 1.50        0.10 0.12 0.16 0.50 0.50     
    WIDTH 4.50        0.10 0.12 0.16 0.50 1.50 ;
    MINENCLOSEDAREA  0.20 ;
    PROPERTY LEF57_MINSTEP "MINSTEP 0.10 MAXEDGES 1 ;" ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    MINIMUMCUT 2 WIDTH 0.30 ;
    MINIMUMCUT 4 WIDTH 0.70 ;
    MINIMUMCUT 2 WIDTH 0.3 LENGTH  0.3 WITHIN 0.8 ;
    MINIMUMCUT 2 WIDTH 2.0 LENGTH  2.0 WITHIN 2 ;
    MINIMUMCUT 2 WIDTH 3.0 LENGTH 10.0 WITHIN 5 ;
    ANTENNACUMAREARATIO 4996 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 4996 ) ( 0.059 4996 ) ( 0.06 43017 ) ( 1 43436 ) ) ;
    THICKNESS 0.22 ;
    HEIGHT 2.62 ;
    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
    FILLACTIVESPACING 0.61 ;
    RESISTANCE RPERSQ       1.4000e-01 ;
    CAPACITANCE CPERSQDIST  3.5957e-04 ;
    EDGECAPACITANCE        10.4751e-05 ;
END M7

LAYER VIA7
    TYPE CUT ;
    SPACING 0.54 ;
    SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;
    ENCLOSURE BELOW 0.08 0.02 ;
    ENCLOSURE ABOVE 0.08 0.02 ;
    ANTENNAAREARATIO 19 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 19 ) ( 0.059 19 ) ( 0.06 903 ) ( 1 1098 ) ) ;
END VIA7

LAYER M8
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    WIDTH 0.40 ;
    MAXWIDTH 12.00 ; 
    PITCH 0.80 ;
    OFFSET 0.40 ;
    AREA 0.565 ;
    SPACINGTABLE
    PARALLELRUNLENGTH 0.00 1.50 4.50     
    WIDTH 0.00        0.40 0.40 0.40     
    WIDTH 1.50        0.40 0.50 0.50      
    WIDTH 4.50        0.40 0.50 1.50 ;
    MINENCLOSEDAREA  0.565 ;
    PROPERTY LEF57_MINSTEP "MINSTEP 0.40 MAXEDGES 1 ;" ;
    MINIMUMCUT 2 WIDTH 1.80 ;
    MINIMUMCUT 2 WIDTH 3.0 LENGTH 10.0 WITHIN 5 ;
    ANTENNACUMAREARATIO 4996 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 4996 ) ( 0.059 4996 ) ( 0.06 50470 ) ( 1 57980 ) ) ;
    THICKNESS 0.9 ;
    HEIGHT 3.435 ;
    MINIMUMDENSITY 20 ;
    MAXIMUMDENSITY 80 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
    FILLACTIVESPACING 1.17 ;
    RESISTANCE RPERSQ       2.2000e-02 ;
    CAPACITANCE CPERSQDIST 10.7397e-05 ;
    EDGECAPACITANCE        15.0247e-05 ;
END M8

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

MAXVIASTACK 4 RANGE M1 M7 ;

VIA VIA1_H DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M1 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA1 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M2 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA1_H

VIA VIA1_V DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M1 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA1 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M2 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA1_V

VIA VIA1_X DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M1 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA1 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M2 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA1_X

VIA VIA1_XR DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M1 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA1 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M2 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA1_XR

VIA VIA2_H DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M2 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA2 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M3 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA2_H

VIA VIA2_V DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M2 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA2 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M3 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA2_V

VIA VIA2_X DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M2 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA2 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M3 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA2_X

VIA VIA2_XR DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M2 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA2 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M3 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA2_XR

VIA VIA3_H DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M3 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA3 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M4 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA3_H

VIA VIA3_V DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M3 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA3 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M4 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA3_V

VIA VIA3_X DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M3 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA3 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M4 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA3_X

VIA VIA3_XR DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M3 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA3 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M4 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA3_XR

VIA VIA4_H DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M4 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA4 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M5 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA4_H

VIA VIA4_V DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M4 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA4 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M5 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA4_V

VIA VIA4_X DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M4 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA4 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M5 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA4_X

VIA VIA4_XR DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M4 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA4 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M5 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA4_XR

VIA VIA5_H DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M5 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA5 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M6 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA5_H

VIA VIA5_V DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M5 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA5 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M6 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA5_V

VIA VIA5_X DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M5 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA5 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M6 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA5_X

VIA VIA5_XR DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M5 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA5 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M6 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA5_XR

VIA VIA6_H DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M6 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA6 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M7 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA6_H

VIA VIA6_V DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M6 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA6 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M7 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA6_V

VIA VIA6_X DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M6 ;
        RECT -0.05 -0.09 0.05 0.09 ;
    LAYER VIA6 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M7 ;
        RECT -0.09 -0.05 0.09 0.05 ;
END VIA6_X

VIA VIA6_XR DEFAULT
    RESISTANCE 1.5000e+00 ;
    LAYER M6 ;
        RECT -0.09 -0.05 0.09 0.05 ;
    LAYER VIA6 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M7 ;
        RECT -0.05 -0.09 0.05 0.09 ;
END VIA6_XR

VIA VIA7_H DEFAULT
    RESISTANCE 2.2000e-01 ;
    LAYER M7 ;
        RECT -0.26 -0.2 0.26 0.2 ;
    LAYER VIA7 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER M8 ;
        RECT -0.26 -0.2 0.26 0.2 ;
END VIA7_H

VIA VIA7_V DEFAULT
    RESISTANCE 2.2000e-01 ;
    LAYER M7 ;
        RECT -0.2 -0.26 0.2 0.26 ;
    LAYER VIA7 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER M8 ;
        RECT -0.2 -0.26 0.2 0.26 ;
END VIA7_V

VIA VIA7_X DEFAULT
    RESISTANCE 2.2000e-01 ;
    LAYER M7 ;
        RECT -0.26 -0.2 0.26 0.2 ;
    LAYER VIA7 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER M8 ;
        RECT -0.2 -0.26 0.2 0.26 ;
END VIA7_X

VIA VIA7_XR DEFAULT
    RESISTANCE 2.2000e-01 ;
    LAYER M7 ;
        RECT -0.2 -0.26 0.2 0.26 ;
    LAYER VIA7 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER M8 ;
        RECT -0.26 -0.2 0.26 0.2 ;
END VIA7_XR

VIA VIA1_2CUT_E DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M1 ;
        RECT -0.09 -0.05 0.29 0.05 ;
    LAYER VIA1 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT 0.15 -0.05 0.25 0.05 ;
    LAYER M2 ;
        RECT -0.09 -0.05 0.29 0.05 ;
END VIA1_2CUT_E

VIA VIA1_2CUT_W DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M1 ;
        RECT -0.29 -0.05 0.09 0.05 ;
    LAYER VIA1 ;
        RECT -0.25 -0.05 -0.15 0.05 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M2 ;
        RECT -0.29 -0.05 0.09 0.05 ;
END VIA1_2CUT_W

VIA VIA1_2CUT_N DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M1 ;
        RECT -0.05 -0.09 0.05 0.29 ;
    LAYER VIA1 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT -0.05 0.15 0.05 0.25 ;
    LAYER M2 ;
        RECT -0.05 -0.09 0.05 0.29 ;
END VIA1_2CUT_N

VIA VIA1_2CUT_S DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M1 ;
        RECT -0.05 -0.29 0.05 0.09 ;
    LAYER VIA1 ;
        RECT -0.05 -0.25 0.05 -0.15 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M2 ;
        RECT -0.05 -0.29 0.05 0.09 ;
END VIA1_2CUT_S

VIA VIA2_2CUT_E DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M2 ;
        RECT -0.09 -0.05 0.29 0.05 ;
    LAYER VIA2 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT 0.15 -0.05 0.25 0.05 ;
    LAYER M3 ;
        RECT -0.09 -0.05 0.29 0.05 ;
END VIA2_2CUT_E

VIA VIA2_2CUT_W DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M2 ;
        RECT -0.29 -0.05 0.09 0.05 ;
    LAYER VIA2 ;
        RECT -0.25 -0.05 -0.15 0.05 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M3 ;
        RECT -0.29 -0.05 0.09 0.05 ;
END VIA2_2CUT_W

VIA VIA2_2CUT_N DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M2 ;
        RECT -0.05 -0.09 0.05 0.29 ;
    LAYER VIA2 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT -0.05 0.15 0.05 0.25 ;
    LAYER M3 ;
        RECT -0.05 -0.09 0.05 0.29 ;
END VIA2_2CUT_N

VIA VIA2_2CUT_S DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M2 ;
        RECT -0.05 -0.29 0.05 0.09 ;
    LAYER VIA2 ;
        RECT -0.05 -0.25 0.05 -0.15 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M3 ;
        RECT -0.05 -0.29 0.05 0.09 ;
END VIA2_2CUT_S

VIA VIA3_2CUT_E DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M3 ;
        RECT -0.09 -0.05 0.29 0.05 ;
    LAYER VIA3 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT 0.15 -0.05 0.25 0.05 ;
    LAYER M4 ;
        RECT -0.09 -0.05 0.29 0.05 ;
END VIA3_2CUT_E

VIA VIA3_2CUT_W DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M3 ;
        RECT -0.29 -0.05 0.09 0.05 ;
    LAYER VIA3 ;
        RECT -0.25 -0.05 -0.15 0.05 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M4 ;
        RECT -0.29 -0.05 0.09 0.05 ;
END VIA3_2CUT_W

VIA VIA3_2CUT_N DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M3 ;
        RECT -0.05 -0.09 0.05 0.29 ;
    LAYER VIA3 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT -0.05 0.15 0.05 0.25 ;
    LAYER M4 ;
        RECT -0.05 -0.09 0.05 0.29 ;
END VIA3_2CUT_N

VIA VIA3_2CUT_S DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M3 ;
        RECT -0.05 -0.29 0.05 0.09 ;
    LAYER VIA3 ;
        RECT -0.05 -0.25 0.05 -0.15 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M4 ;
        RECT -0.05 -0.29 0.05 0.09 ;
END VIA3_2CUT_S

VIA VIA4_2CUT_E DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M4 ;
        RECT -0.09 -0.05 0.29 0.05 ;
    LAYER VIA4 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT 0.15 -0.05 0.25 0.05 ;
    LAYER M5 ;
        RECT -0.09 -0.05 0.29 0.05 ;
END VIA4_2CUT_E

VIA VIA4_2CUT_W DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M4 ;
        RECT -0.29 -0.05 0.09 0.05 ;
    LAYER VIA4 ;
        RECT -0.25 -0.05 -0.15 0.05 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M5 ;
        RECT -0.29 -0.05 0.09 0.05 ;
END VIA4_2CUT_W

VIA VIA4_2CUT_N DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M4 ;
        RECT -0.05 -0.09 0.05 0.29 ;
    LAYER VIA4 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT -0.05 0.15 0.05 0.25 ;
    LAYER M5 ;
        RECT -0.05 -0.09 0.05 0.29 ;
END VIA4_2CUT_N

VIA VIA4_2CUT_S DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M4 ;
        RECT -0.05 -0.29 0.05 0.09 ;
    LAYER VIA4 ;
        RECT -0.05 -0.25 0.05 -0.15 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M5 ;
        RECT -0.05 -0.29 0.05 0.09 ;
END VIA4_2CUT_S

VIA VIA5_2CUT_E DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M5 ;
        RECT -0.09 -0.05 0.29 0.05 ;
    LAYER VIA5 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT 0.15 -0.05 0.25 0.05 ;
    LAYER M6 ;
        RECT -0.09 -0.05 0.29 0.05 ;
END VIA5_2CUT_E

VIA VIA5_2CUT_W DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M5 ;
        RECT -0.29 -0.05 0.09 0.05 ;
    LAYER VIA5 ;
        RECT -0.25 -0.05 -0.15 0.05 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M6 ;
        RECT -0.29 -0.05 0.09 0.05 ;
END VIA5_2CUT_W

VIA VIA5_2CUT_N DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M5 ;
        RECT -0.05 -0.09 0.05 0.29 ;
    LAYER VIA5 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT -0.05 0.15 0.05 0.25 ;
    LAYER M6 ;
        RECT -0.05 -0.09 0.05 0.29 ;
END VIA5_2CUT_N

VIA VIA5_2CUT_S DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M5 ;
        RECT -0.05 -0.29 0.05 0.09 ;
    LAYER VIA5 ;
        RECT -0.05 -0.25 0.05 -0.15 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M6 ;
        RECT -0.05 -0.29 0.05 0.09 ;
END VIA5_2CUT_S

VIA VIA6_2CUT_E DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M6 ;
        RECT -0.09 -0.05 0.29 0.05 ;
    LAYER VIA6 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT 0.15 -0.05 0.25 0.05 ;
    LAYER M7 ;
        RECT -0.09 -0.05 0.29 0.05 ;
END VIA6_2CUT_E

VIA VIA6_2CUT_W DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M6 ;
        RECT -0.29 -0.05 0.09 0.05 ;
    LAYER VIA6 ;
        RECT -0.25 -0.05 -0.15 0.05 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M7 ;
        RECT -0.29 -0.05 0.09 0.05 ;
END VIA6_2CUT_W

VIA VIA6_2CUT_N DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M6 ;
        RECT -0.05 -0.09 0.05 0.29 ;
    LAYER VIA6 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        RECT -0.05 0.15 0.05 0.25 ;
    LAYER M7 ;
        RECT -0.05 -0.09 0.05 0.29 ;
END VIA6_2CUT_N

VIA VIA6_2CUT_S DEFAULT
    RESISTANCE 7.5000e-01 ;
    LAYER M6 ;
        RECT -0.05 -0.29 0.05 0.09 ;
    LAYER VIA6 ;
        RECT -0.05 -0.25 0.05 -0.15 ;
        RECT -0.05 -0.05 0.05 0.05 ;
    LAYER M7 ;
        RECT -0.05 -0.29 0.05 0.09 ;
END VIA6_2CUT_S

VIA VIA7_2CUT_E DEFAULT
    RESISTANCE 1.1000e-01 ;
    LAYER M7 ;
        RECT -0.26 -0.2 0.96 0.2 ;
    LAYER VIA7 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        RECT 0.52 -0.18 0.88 0.18 ;
    LAYER M8 ;
        RECT -0.26 -0.2 0.96 0.2 ;
END VIA7_2CUT_E

VIA VIA7_2CUT_W DEFAULT
    RESISTANCE 1.1000e-01 ;
    LAYER M7 ;
        RECT -0.96 -0.2 0.26 0.2 ;
    LAYER VIA7 ;
        RECT -0.88 -0.18 -0.52 0.18 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER M8 ;
        RECT -0.96 -0.2 0.26 0.2 ;
END VIA7_2CUT_W

VIA VIA7_2CUT_N DEFAULT
    RESISTANCE 1.1000e-01 ;
    LAYER M7 ;
        RECT -0.2 -0.26 0.2 0.96 ;
    LAYER VIA7 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        RECT -0.18 0.52 0.18 0.88 ;
    LAYER M8 ;
        RECT -0.2 -0.26 0.2 0.96 ;
END VIA7_2CUT_N

VIA VIA7_2CUT_S DEFAULT
    RESISTANCE 1.1000e-01 ;
    LAYER M7 ;
        RECT -0.2 -0.96 0.2 0.26 ;
    LAYER VIA7 ;
        RECT -0.18 -0.88 0.18 -0.52 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER M8 ;
        RECT -0.2 -0.96 0.2 0.26 ;
END VIA7_2CUT_S

VIA VIA1_4CUT DEFAULT
    RESISTANCE 3.75e-01 ;
    LAYER M1 ;
        RECT -0.165 -0.205 0.165 0.205 ;
    LAYER VIA1 ;
        RECT -0.165 -0.165 -0.065 -0.065 ;
        RECT 0.065 -0.165 0.165 -0.065 ;
        RECT -0.165 0.065 -0.065 0.165 ;
        RECT 0.065 0.065 0.165 0.165 ;
    LAYER M2 ;
        RECT -0.205 -0.165 0.205 0.165 ;
END VIA1_4CUT

VIA VIA2_4CUT DEFAULT
    RESISTANCE 3.75e-01 ;
    LAYER M2 ;
        RECT -0.205 -0.165 0.205 0.165 ;
    LAYER VIA2 ;
        RECT -0.165 -0.165 -0.065 -0.065 ;
        RECT 0.065 -0.165 0.165 -0.065 ;
        RECT -0.165 0.065 -0.065 0.165 ;
        RECT 0.065 0.065 0.165 0.165 ;
    LAYER M3 ;
        RECT -0.205 -0.165 0.205 0.165 ;
END VIA2_4CUT

VIA VIA3_4CUT DEFAULT
    RESISTANCE 3.75e-01 ;
    LAYER M3 ;
        RECT -0.205 -0.165 0.205 0.165 ;
    LAYER VIA3 ;
        RECT -0.165 -0.165 -0.065 -0.065 ;
        RECT 0.065 -0.165 0.165 -0.065 ;
        RECT -0.165 0.065 -0.065 0.165 ;
        RECT 0.065 0.065 0.165 0.165 ;
    LAYER M4 ;
        RECT -0.205 -0.165 0.205 0.165 ;
END VIA3_4CUT

VIA VIA4_4CUT DEFAULT
    RESISTANCE 3.75e-01 ;
    LAYER M4 ;
        RECT -0.205 -0.165 0.205 0.165 ;
    LAYER VIA4 ;
        RECT -0.165 -0.165 -0.065 -0.065 ;
        RECT 0.065 -0.165 0.165 -0.065 ;
        RECT -0.165 0.065 -0.065 0.165 ;
        RECT 0.065 0.065 0.165 0.165 ;
    LAYER M5 ;
        RECT -0.205 -0.165 0.205 0.165 ;
END VIA4_4CUT

VIA VIA5_4CUT DEFAULT
    RESISTANCE 3.75e-01 ;
    LAYER M5 ;
        RECT -0.205 -0.165 0.205 0.165 ;
    LAYER VIA5 ;
        RECT -0.165 -0.165 -0.065 -0.065 ;
        RECT 0.065 -0.165 0.165 -0.065 ;
        RECT -0.165 0.065 -0.065 0.165 ;
        RECT 0.065 0.065 0.165 0.165 ;
    LAYER M6 ;
        RECT -0.205 -0.165 0.205 0.165 ;
END VIA5_4CUT

VIA VIA6_4CUT DEFAULT
    RESISTANCE 3.75e-01 ;
    LAYER M6 ;
        RECT -0.205 -0.165 0.205 0.165 ;
    LAYER VIA6 ;
        RECT -0.165 -0.165 -0.065 -0.065 ;
        RECT 0.065 -0.165 0.165 -0.065 ;
        RECT -0.165 0.065 -0.065 0.165 ;
        RECT 0.065 0.065 0.165 0.165 ;
    LAYER M7 ;
        RECT -0.205 -0.165 0.205 0.165 ;
END VIA6_4CUT

VIA VIA7_4CUT DEFAULT
    RESISTANCE 5.50e-02 ;
    LAYER M7 ;
        RECT -0.71 -0.65 0.71 0.65 ;
    LAYER VIA7 ;
        RECT -0.63 -0.63 -0.27 -0.27 ;
        RECT 0.27 -0.63 0.63 -0.27 ;
        RECT -0.63 0.27 -0.27 0.63 ;
        RECT 0.27 0.27 0.63 0.63 ;
    LAYER M8 ;
        RECT -0.71 -0.65 0.71 0.65 ;
END VIA7_4CUT

VIARULE via1Array GENERATE
    LAYER M1 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER M2 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER VIA1 ;
        RECT -0.050 -0.050 0.050 0.050 ;
        SPACING 0.23 BY 0.23 ;
END via1Array

VIARULE via2Array GENERATE
    LAYER M2 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER M3 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER VIA2 ;
        RECT -0.050 -0.050 0.050 0.050 ;
        SPACING 0.23 BY 0.23 ;
END via2Array

VIARULE via3Array GENERATE
    LAYER M3 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER M4 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER VIA3 ;
        RECT -0.050 -0.050 0.050 0.050 ;
        SPACING 0.23 BY 0.23 ;
END via3Array

VIARULE via4Array GENERATE
    LAYER M4 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER M5 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER VIA4 ;
        RECT -0.050 -0.050 0.050 0.050 ;
        SPACING 0.23 BY 0.23 ;
END via4Array

VIARULE via5Array GENERATE
    LAYER M5 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER M6 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER VIA5 ;
        RECT -0.050 -0.050 0.050 0.050 ;
        SPACING 0.23 BY 0.23 ;
END via5Array

VIARULE via6Array GENERATE
    LAYER M6 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER M7 ;
        ENCLOSURE 0.04 0.0 ;

    LAYER VIA6 ;
        RECT -0.050 -0.050 0.050 0.050 ;
        SPACING 0.23 BY 0.23 ;
END via6Array

VIARULE via7Array GENERATE
    LAYER M7 ;
        ENCLOSURE 0.08 0.02 ;

    LAYER M8 ;
        ENCLOSURE 0.08 0.02 ;

    LAYER VIA7 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        SPACING 0.90 BY 0.90 ;
END via7Array


VIARULE TURNM1 GENERATE
    LAYER M1 ;
        DIRECTION vertical ;

    LAYER M1 ;
        DIRECTION horizontal ;
END TURNM1

VIARULE TURNM2 GENERATE
    LAYER M2 ;
        DIRECTION vertical ;
        
    LAYER M2 ;
        DIRECTION horizontal ;
END TURNM2
    
VIARULE TURNM3 GENERATE
    LAYER M3 ;
        DIRECTION vertical ;

    LAYER M3 ;
        DIRECTION horizontal ;
END TURNM3

VIARULE TURNM4 GENERATE
    LAYER M4 ;
        DIRECTION vertical ;

    LAYER M4 ;
        DIRECTION horizontal ;
END TURNM4

VIARULE TURNM5 GENERATE
    LAYER M5 ;
        DIRECTION vertical ;

    LAYER M5 ;
        DIRECTION horizontal ;
END TURNM5

VIARULE TURNM6 GENERATE
    LAYER M6 ;
        DIRECTION vertical ;

    LAYER M6 ;
        DIRECTION horizontal ;
END TURNM6

VIARULE TURNM7 GENERATE
    LAYER M7 ;
        DIRECTION vertical ;

    LAYER M7 ;
        DIRECTION horizontal ;
END TURNM7

VIARULE TURNM8 GENERATE
    LAYER M8 ;
        DIRECTION vertical ;

    LAYER M8 ;
        DIRECTION horizontal ;
END TURNM8

# Updated by Maxx Seminario for higher DRC Compliance of Innovus for Myshkin chip

SPACING 
    SAMENET M1 M1 0.09  ; 
    SAMENET M2 M2 0.13 STACK ;
    SAMENET M3 M3 0.13 STACK ;
    SAMENET M4 M4 0.13 STACK ;
    SAMENET M5 M5 0.13 STACK ;
    SAMENET M6 M6 0.13 STACK ;
    SAMENET M7 M7 0.13 STACK ;
    SAMENET M8 M8 0.40  ;
    SAMENET VIA1 VIA1 0.10  ;
    SAMENET VIA2 VIA2 0.10  ;
    SAMENET VIA3 VIA3 0.10  ;
    SAMENET VIA4 VIA4 0.10  ;
    SAMENET VIA5 VIA5 0.10  ;
    SAMENET VIA6 VIA6 0.10  ;
    SAMENET VIA7 VIA7 0.34  ;
    SAMENET VIA1 VIA2 0.0 STACK ;
    SAMENET VIA2 VIA3 0.0 STACK ;
    SAMENET VIA3 VIA4 0.0 STACK ;
    SAMENET VIA4 VIA5 0.0 STACK ;
    SAMENET VIA5 VIA6 0.0 STACK ;
    SAMENET VIA6 VIA7 0.0 STACK ;
END SPACING

END LIBRARY
