

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO MCU 
  PIN resetn_in 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 25.762 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 113.397 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 974.013 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4292.32 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6 ;
  END resetn_in
  PIN resetn_out 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.474 LAYER M2 ;
  END resetn_out
  PIN resetn_dir 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6654 LAYER M2 ;
  END resetn_dir
  PIN resetn_ren 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1086 LAYER M2 ;
  END resetn_ren
  PIN prt1_in[7] 
    ANTENNAPARTIALMETALAREA 4.0155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6682 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.358 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.2192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 292.317 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1270.5 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt1_in[7]
  PIN prt1_in[6] 
    ANTENNAPARTIALMETALAREA 23.4525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 103.191 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.626 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.9984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 137.023 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 601.503 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.734684 LAYER VIA3 ;
  END prt1_in[6]
  PIN prt1_in[5] 
    ANTENNAPARTIALMETALAREA 1.5525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.831 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.714 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.6736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2577 LAYER M3 ; 
    ANTENNAMAXAREACAR 249.791 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1100.06 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.786164 LAYER VIA3 ;
  END prt1_in[5]
  PIN prt1_in[4] 
    ANTENNAPARTIALMETALAREA 1.7525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.711 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.95 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1305 LAYER M3 ; 
    ANTENNAMAXAREACAR 138.076 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 607.304 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 1.09665 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.638 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8512 LAYER M4 ;
    ANTENNAGATEAREA 0.1305 LAYER M4 ; 
    ANTENNAMAXAREACAR 142.965 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 629.153 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 1.24991 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.282 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4848 LAYER M5 ;
    ANTENNAGATEAREA 0.2577 LAYER M5 ; 
    ANTENNAMAXAREACAR 155.701 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 685.361 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.24991 LAYER VIA5 ;
  END prt1_in[4]
  PIN prt1_in[3] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5142 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.968 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 LAYER M4 ; 
    ANTENNAMAXAREACAR 27.3687 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 38.6211 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.707547 LAYER VIA4 ;
  END prt1_in[3]
  PIN prt1_in[2] 
    ANTENNAPARTIALMETALAREA 4.5935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.2554 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.378 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.7072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0595 LAYER M3 ; 
    ANTENNAMAXAREACAR 260.039 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1145.03 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.672269 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.346 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3664 LAYER M4 ;
    ANTENNAGATEAREA 0.1633 LAYER M4 ; 
    ANTENNAMAXAREACAR 274.405 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1208.51 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.672269 LAYER VIA4 ;
  END prt1_in[2]
  PIN prt1_in[1] 
    ANTENNAPARTIALMETALAREA 1.2935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.566 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.3344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 165.127 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 726.304 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.339751 LAYER VIA3 ;
  END prt1_in[1]
  PIN prt1_in[0] 
    ANTENNAPARTIALMETALAREA 24.8355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 109.276 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.1568 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M3 ; 
    ANTENNAMAXAREACAR 570.598 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2508.59 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.63265 LAYER VIA3 ;
  END prt1_in[0]
  PIN prt1_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.834 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.3136 LAYER M2 ;
  END prt1_out[7]
  PIN prt1_out[6] 
    ANTENNAPARTIALMETALAREA 0.816 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5904 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.586 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0224 LAYER M3 ;
  END prt1_out[6]
  PIN prt1_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[5]
  PIN prt1_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[4]
  PIN prt1_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[3]
  PIN prt1_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[2]
  PIN prt1_out[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[1]
  PIN prt1_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.495 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.666 LAYER M2 ;
  END prt1_out[0]
  PIN prt1_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.5795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8378 LAYER M2 ;
  END prt1_dir[7]
  PIN prt1_dir[6] 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3046 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4784 LAYER M3 ;
  END prt1_dir[6]
  PIN prt1_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
  END prt1_dir[5]
  PIN prt1_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
  END prt1_dir[4]
  PIN prt1_dir[3] 
    ANTENNAPARTIALMETALAREA 0.3565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5686 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.686 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.0624 LAYER M3 ;
  END prt1_dir[3]
  PIN prt1_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
  END prt1_dir[2]
  PIN prt1_dir[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[1]
  PIN prt1_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.1945 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 53.7438 LAYER M2 ;
  END prt1_dir[0]
  PIN prt1_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5082 LAYER M2 ;
  END prt1_ren[7]
  PIN prt1_ren[6] 
    ANTENNAPARTIALMETALAREA 1.2005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2822 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.686 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4624 LAYER M3 ;
  END prt1_ren[6]
  PIN prt1_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.5875 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.273 LAYER M2 ;
  END prt1_ren[5]
  PIN prt1_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2 ;
  END prt1_ren[4]
  PIN prt1_ren[3] 
    ANTENNAPARTIALMETALAREA 0.2275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.001 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9488 LAYER M3 ;
  END prt1_ren[3]
  PIN prt1_ren[2] 
    ANTENNAPARTIALMETALAREA 1.5455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.612 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9808 LAYER M3 ;
  END prt1_ren[2]
  PIN prt1_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.3705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 54.5182 LAYER M2 ;
  END prt1_ren[1]
  PIN prt1_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.7305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.1022 LAYER M2 ;
  END prt1_ren[0]
  PIN prt2_in[7] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 26.046 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 114.646 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M6 ; 
    ANTENNAMAXAREACAR 766.274 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3366.55 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.88184 LAYER VIA6 ;
  END prt2_in[7]
  PIN prt2_in[6] 
    ANTENNAPARTIALMETALAREA 0.7175 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.201 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 33.4438 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 142.409 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END prt2_in[6]
  PIN prt2_in[5] 
    ANTENNAPARTIALMETALAREA 0.6755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9722 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.78796 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 29.187 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0925926 LAYER VIA2 ;
  END prt2_in[5]
  PIN prt2_in[4] 
    ANTENNAPARTIALMETALAREA 0.5955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6202 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.626 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.7984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 169.308 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 744.386 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt2_in[4]
  PIN prt2_in[3] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3916 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.432 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M4 ; 
    ANTENNAMAXAREACAR 16.8145 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 23.1195 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.314465 LAYER VIA4 ;
  END prt2_in[3]
  PIN prt2_in[2] 
    ANTENNAPARTIALMETALAREA 0.5395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3738 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.29245 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 13.9979 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.104822 LAYER VIA2 ;
  END prt2_in[2]
  PIN prt2_in[1] 
    ANTENNAPARTIALMETALAREA 0.3555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5642 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 26.266 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 115.614 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0595 LAYER M3 ; 
    ANTENNAMAXAREACAR 474.87 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2079.55 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.672269 LAYER VIA3 ;
  END prt2_in[1]
  PIN prt2_in[0] 
    ANTENNAPARTIALMETALAREA 0.5535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4794 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.246 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.5264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M3 ; 
    ANTENNAMAXAREACAR 86.3684 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 378.186 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.209644 LAYER VIA3 ;
  END prt2_in[0]
  PIN prt2_out[7] 
    ANTENNAPARTIALMETALAREA 0.691 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.9168 LAYER M3 ;
  END prt2_out[7]
  PIN prt2_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.681 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0404 LAYER M2 ;
  END prt2_out[6]
  PIN prt2_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.777 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5508 LAYER M2 ;
  END prt2_out[5]
  PIN prt2_out[4] 
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.4368 LAYER M3 ;
  END prt2_out[4]
  PIN prt2_out[3] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.914 LAYER M2 ;
  END prt2_out[3]
  PIN prt2_out[2] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.266 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.8144 LAYER M3 ;
  END prt2_out[2]
  PIN prt2_out[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.459 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0196 LAYER M2 ;
  END prt2_out[1]
  PIN prt2_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.292 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M2 ;
  END prt2_out[0]
  PIN prt2_dir[7] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2254 LAYER M2 ;
  END prt2_dir[7]
  PIN prt2_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7015 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1306 LAYER M2 ;
  END prt2_dir[6]
  PIN prt2_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3198 LAYER M2 ;
  END prt2_dir[5]
  PIN prt2_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2 ;
  END prt2_dir[4]
  PIN prt2_dir[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3706 LAYER M2 ;
  END prt2_dir[3]
  PIN prt2_dir[2] 
    ANTENNAPARTIALMETALAREA 0.431 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8964 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.978 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.9472 LAYER M3 ;
  END prt2_dir[2]
  PIN prt2_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3046 LAYER M2 ;
  END prt2_dir[1]
  PIN prt2_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2506 LAYER M2 ;
  END prt2_dir[0]
  PIN prt2_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4102 LAYER M2 ;
  END prt2_ren[7]
  PIN prt2_ren[6] 
    ANTENNAPARTIALMETALAREA 0.6205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7302 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.706 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5504 LAYER M3 ;
  END prt2_ren[6]
  PIN prt2_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2362 LAYER M2 ;
  END prt2_ren[5]
  PIN prt2_ren[4] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.518 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.7232 LAYER M3 ;
  END prt2_ren[4]
  PIN prt2_ren[3] 
    ANTENNAPARTIALMETALAREA 0.6075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.673 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8544 LAYER M3 ;
  END prt2_ren[3]
  PIN prt2_ren[2] 
    ANTENNAPARTIALMETALAREA 0.647 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8468 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.3855 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5402 LAYER M3 ;
  END prt2_ren[2]
  PIN prt2_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4794 LAYER M2 ;
  END prt2_ren[1]
  PIN prt2_ren[0] 
    ANTENNAPARTIALMETALAREA 0.4675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.057 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.266 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.6144 LAYER M3 ;
  END prt2_ren[0]
  PIN prt3_in[7] 
    ANTENNAPARTIALMETALAREA 18.1685 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 80.0294 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 672.039 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2958.76 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2 ;
  END prt3_in[7]
  PIN prt3_in[6] 
    ANTENNAPARTIALMETALAREA 9.5105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 41.8902 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 352.555 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 1551.41 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2 ;
  END prt3_in[6]
  PIN prt3_in[5] 
    ANTENNAPARTIALMETALAREA 6.8725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.239 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 14.464 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.7296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M3 ; 
    ANTENNAMAXAREACAR 408.863 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1790.57 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 2.71003 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.498 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6352 LAYER M4 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 423.295 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1854.49 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.71003 LAYER VIA4 ;
  END prt3_in[5]
  PIN prt3_in[4] 
    ANTENNAPARTIALMETALAREA 0.4395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9338 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.006 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.0704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 152.263 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 671.113 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3 ;
  END prt3_in[4]
  PIN prt3_in[3] 
    ANTENNAPARTIALMETALAREA 1.1955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2602 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.068 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.3872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M3 ; 
    ANTENNAMAXAREACAR 538.103 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2370.77 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 1.89702 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4032 LAYER M4 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 549.837 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 2422.82 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 2.0897 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 8.126 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 35.7984 LAYER M5 ;
    ANTENNAGATEAREA 0.1707 LAYER M5 ; 
    ANTENNAMAXAREACAR 597.441 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2632.54 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.0897 LAYER VIA5 ;
  END prt3_in[3]
  PIN prt3_in[2] 
    ANTENNAPARTIALMETALAREA 0.5755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 481.688 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2126.09 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3 ;
  END prt3_in[2]
  PIN prt3_in[1] 
    ANTENNAPARTIALMETALAREA 14.9555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.8042 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.338 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.1312 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 189.756 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 814.465 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[1]
  PIN prt3_in[0] 
    ANTENNAPARTIALMETALAREA 1.8525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.151 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.5568 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 301.078 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1309.04 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt3_in[0]
  PIN prt3_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.801 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.1684 LAYER M2 ;
  END prt3_out[7]
  PIN prt3_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.339 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9796 LAYER M2 ;
  END prt3_out[6]
  PIN prt3_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.137 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6468 LAYER M2 ;
  END prt3_out[5]
  PIN prt3_out[4] 
    ANTENNAPARTIALMETALAREA 0.316 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.4448 LAYER M3 ;
  END prt3_out[4]
  PIN prt3_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.137 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6468 LAYER M2 ;
  END prt3_out[3]
  PIN prt3_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 10.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 45.848 LAYER M2 ;
  END prt3_out[2]
  PIN prt3_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.378 LAYER M2 ;
  END prt3_out[1]
  PIN prt3_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.901 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2084 LAYER M2 ;
  END prt3_out[0]
  PIN prt3_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.8395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 60.9818 LAYER M2 ;
  END prt3_dir[7]
  PIN prt3_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 7.5615 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.3146 LAYER M2 ;
  END prt3_dir[6]
  PIN prt3_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt3_dir[5]
  PIN prt3_dir[4] 
    ANTENNAPARTIALMETALAREA 0.2565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.902 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 52.4128 LAYER M3 ;
  END prt3_dir[4]
  PIN prt3_dir[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt3_dir[3]
  PIN prt3_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.2545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.2078 LAYER M2 ;
  END prt3_dir[2]
  PIN prt3_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.9765 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.6286 LAYER M2 ;
  END prt3_dir[1]
  PIN prt3_dir[0] 
    ANTENNAPARTIALMETALAREA 2.8695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.3728 LAYER M3 ;
  END prt3_dir[0]
  PIN prt3_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.3675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.905 LAYER M2 ;
  END prt3_ren[7]
  PIN prt3_ren[6] 
    ANTENNAPARTIALMETALAREA 4.7385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.8934 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4928 LAYER M3 ;
  END prt3_ren[6]
  PIN prt3_ren[5] 
    ANTENNAPARTIALMETALAREA 4.1005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.0422 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.6368 LAYER M3 ;
  END prt3_ren[5]
  PIN prt3_ren[4] 
    ANTENNAPARTIALMETALAREA 0.3005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.6528 LAYER M3 ;
  END prt3_ren[4]
  PIN prt3_ren[3] 
    ANTENNAPARTIALMETALAREA 1.1855 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2602 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.706 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.1504 LAYER M3 ;
  END prt3_ren[3]
  PIN prt3_ren[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 7.1125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.427 LAYER M2 ;
  END prt3_ren[2]
  PIN prt3_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.3125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 63.107 LAYER M2 ;
  END prt3_ren[1]
  PIN prt3_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.5255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2442 LAYER M2 ;
  END prt3_ren[0]
  PIN prt4_in[7] 
    ANTENNAPARTIALMETALAREA 1.3555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9642 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 26.284 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 115.738 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 258.354 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1136.84 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3 ;
  END prt4_in[7]
  PIN prt4_in[6] 
    ANTENNAPARTIALMETALAREA 2.0355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9562 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.668 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.4272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M3 ; 
    ANTENNAMAXAREACAR 591.237 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2593.78 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 2.71003 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.658 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9392 LAYER M4 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 597.576 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 2622.09 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.71003 LAYER VIA4 ;
  END prt4_in[6]
  PIN prt4_in[5] 
    ANTENNAPARTIALMETALAREA 1.2585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5374 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.794 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.2256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 215.872 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 951.841 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA3 ;
  END prt4_in[5]
  PIN prt4_in[4] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.638 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8512 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 7.518 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.1232 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 98.2719 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 433.74 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA4 ;
  END prt4_in[4]
  PIN prt4_in[3] 
    ANTENNAPARTIALMETALAREA 7.4285 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.7734 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M2 ; 
    ANTENNAMAXAREACAR 74.5371 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 327.346 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.542005 LAYER VIA2 ;
  END prt4_in[3]
  PIN prt4_in[2] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.888 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.7952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 280.955 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1236.58 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
  END prt4_in[2]
  PIN prt4_in[1] 
    ANTENNAPARTIALMETALAREA 7.8905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.7622 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M2 ; 
    ANTENNAMAXAREACAR 215.081 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 947.089 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 217.027 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 956.076 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3 ;
  END prt4_in[1]
  PIN prt4_in[0] 
    ANTENNAPARTIALMETALAREA 0.2925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.287 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 29.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 130.997 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 1107.99 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4862.64 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt4_in[0]
  PIN prt4_out[7] 
    ANTENNAPARTIALMETALAREA 9.292 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.2806 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 65.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 72.512 LAYER M3 ;
  END prt4_out[7]
  PIN prt4_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 10.81 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.9504 LAYER M2 ;
  END prt4_out[6]
  PIN prt4_out[5] 
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.642 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.2822 LAYER M3 ;
  END prt4_out[5]
  PIN prt4_out[4] 
    ANTENNAPARTIALMETALAREA 23.948 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.4022 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.882 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1462 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.162 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3062 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.552 LAYER M5 ;
  END prt4_out[4]
  PIN prt4_out[3] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.998 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.4352 LAYER M3 ;
  END prt4_out[3]
  PIN prt4_out[2] 
    ANTENNAPARTIALMETALAREA 0.499 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1956 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.9024 LAYER M3 ;
  END prt4_out[2]
  PIN prt4_out[1] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[1]
  PIN prt4_out[0] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[0]
  PIN prt4_dir[7] 
    ANTENNAPARTIALMETALAREA 0.3515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5466 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.586 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.0224 LAYER M3 ;
  END prt4_dir[7]
  PIN prt4_dir[6] 
    ANTENNAPARTIALMETALAREA 0.5115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2506 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.886 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.1424 LAYER M3 ;
  END prt4_dir[6]
  PIN prt4_dir[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3222 LAYER M2 ;
  END prt4_dir[5]
  PIN prt4_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.6915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4426 LAYER M2 ;
  END prt4_dir[4]
  PIN prt4_dir[3] 
    ANTENNAPARTIALMETALAREA 0.871 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.998 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.0352 LAYER M3 ;
  END prt4_dir[3]
  PIN prt4_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3418 LAYER M2 ;
  END prt4_dir[2]
  PIN prt4_dir[1] 
    ANTENNAPARTIALMETALAREA 0.5365 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3606 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.218 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 71.4032 LAYER M6 ;
  END prt4_dir[1]
  PIN prt4_dir[0] 
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6 ;
  END prt4_dir[0]
  PIN prt4_ren[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3095 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4058 LAYER M2 ;
  END prt4_ren[7]
  PIN prt4_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.9475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.257 LAYER M2 ;
  END prt4_ren[6]
  PIN prt4_ren[5] 
    ANTENNAPARTIALMETALAREA 1.1105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8862 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.266 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.2144 LAYER M3 ;
  END prt4_ren[5]
  PIN prt4_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.6505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0622 LAYER M2 ;
  END prt4_ren[4]
  PIN prt4_ren[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.5385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0134 LAYER M2 ;
  END prt4_ren[3]
  PIN prt4_ren[2] 
    ANTENNAPARTIALMETALAREA 0.6835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0074 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.5728 LAYER M3 ;
  END prt4_ren[2]
  PIN prt4_ren[1] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_ren[1]
  PIN prt4_ren[0] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.762 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.7968 LAYER M6 ;
  END prt4_ren[0]
  PIN use_dac_glb_bias 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.638 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8512 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.018 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.7232 LAYER M6 ;
  END use_dac_glb_bias
  PIN en_bias_buf 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.498 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.4352 LAYER M4 ;
  END en_bias_buf
  PIN en_bias_gen 
    ANTENNAPARTIALMETALAREA 0.73 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.212 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.882 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.3248 LAYER M4 ;
  END en_bias_gen
  PIN BIAS_ADJ[5] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.842 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.118 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.1632 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.682 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 42.7328 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 196.288 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 862.612 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.678 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0272 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.526 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7584 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.858 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 25.8192 LAYER M6 ;
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3888 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.558 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6992 LAYER M6 ;
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.858 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 30.2192 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 195.867 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 864.903 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA4 ;
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.598 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0752 LAYER M3 ;
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.14 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.304 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 0.366 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M7 ; 
    ANTENNAMAXAREACAR 57.8175 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 256.367 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.7316 LAYER VIA7 ;
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.002 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.8528 LAYER M4 ;
  END BIAS_DBP[13]
  PIN BIAS_DBP[12] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.358 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M3 ;
  END BIAS_DBP[12]
  PIN BIAS_DBP[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.491 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2044 LAYER M2 ;
  END BIAS_DBP[11]
  PIN BIAS_DBP[10] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1562 LAYER M2 ;
  END BIAS_DBP[10]
  PIN BIAS_DBP[9] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
  END BIAS_DBP[9]
  PIN BIAS_DBP[8] 
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3 ;
  END BIAS_DBP[8]
  PIN BIAS_DBP[7] 
    ANTENNAPARTIALMETALAREA 0.127 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5588 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.806 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.0072 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.628 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0512 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.458 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 24.0592 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 338.227 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1491.18 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_DBP[7]
  PIN BIAS_DBP[6] 
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.582 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.338 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7312 LAYER M4 ;
  END BIAS_DBP[6]
  PIN BIAS_DBP[5] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.784 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9376 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.358 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.4192 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.186 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.918 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.6832 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 1.802 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9728 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M7 ; 
    ANTENNAMAXAREACAR 113.883 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 504.704 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.5873 LAYER VIA7 ;
  END BIAS_DBP[5]
  PIN BIAS_DBP[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
  END BIAS_DBP[4]
  PIN BIAS_DBP[3] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.7664 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5152 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.446 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4064 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.458 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 28.4592 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 2.942 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9888 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 226.689 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 1001.28 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA7 ;
  END BIAS_DBP[3]
  PIN BIAS_DBP[2] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.0676 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 12.806 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 56.3904 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 637.181 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2809.09 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_DBP[2]
  PIN BIAS_DBP[1] 
    ANTENNAPARTIALMETALAREA 0.199 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9196 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.546 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8464 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.698 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5592 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.002 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4528 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.924 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7536 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 102.325 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 453.847 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA6 ;
  END BIAS_DBP[1]
  PIN BIAS_DBP[0] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.5635 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9234 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.298 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.1552 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.526 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7584 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.6 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 20.328 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 107.337 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 476.123 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6 ;
  END BIAS_DBP[0]
  PIN BIAS_DBN[13] 
    ANTENNAPARTIALMETALAREA 0.408 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7952 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.398 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.9952 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.322 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0608 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.036 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.8464 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 152.333 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 668.277 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_DBN[13]
  PIN BIAS_DBN[12] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.318 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4432 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.222 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.6208 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.616 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 37.9984 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 233.532 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1030.77 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA6 ;
  END BIAS_DBN[12]
  PIN BIAS_DBN[11] 
    ANTENNAPARTIALMETALAREA 0.031 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.786 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.142 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6688 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.378 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 36.9072 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 288.683 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1274.06 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_DBN[11]
  PIN BIAS_DBN[10] 
    ANTENNAPARTIALMETALAREA 0.4895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1978 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.768 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.8672 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 5.238 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0912 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.266 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 2.418 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 10.6832 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 121.908 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 538.753 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_DBN[10]
  PIN BIAS_DBN[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.934 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0416 LAYER M2 ;
  END BIAS_DBN[9]
  PIN BIAS_DBN[8] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.146 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M3 ;
  END BIAS_DBN[8]
  PIN BIAS_DBN[7] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.389 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7556 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.9584 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.958 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.4592 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 114.917 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 509.483 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_DBN[7]
  PIN BIAS_DBN[6] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.826 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6784 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.206 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.5504 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.278 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 36.4672 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 240.65 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1061.98 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_DBN[6]
  PIN BIAS_DBN[5] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.802 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 43.1728 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 231.756 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1022.53 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA6 ;
  END BIAS_DBN[5]
  PIN BIAS_DBN[4] 
    ANTENNAPARTIALMETALAREA 0.0295 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.702 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.9328 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.658 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 42.5392 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER M6 ; 
    ANTENNAMAXAREACAR 256.872 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1132.81 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.4245 LAYER VIA6 ;
  END BIAS_DBN[4]
  PIN BIAS_DBN[3] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.738 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6912 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.086 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4224 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.978 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 30.7472 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 124.874 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 551.403 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_DBN[3]
  PIN BIAS_DBN[2] 
    ANTENNAPARTIALMETALAREA 0.8785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9094 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 9.388 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.3952 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.762 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1968 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 54.4745 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 241.44 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA5 ;
  END BIAS_DBN[2]
  PIN BIAS_DBN[1] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.488 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.4352 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.1632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.278 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 18.8672 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 185.51 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 817.984 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6 ;
  END BIAS_DBN[1]
  PIN BIAS_DBN[0] 
    ANTENNAPARTIALMETALAREA 0.0315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1386 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.1328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 10.862 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 47.8368 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.338 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3312 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 120.508 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 533.126 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA5 ;
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.063 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3212 LAYER M2 ;
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12] 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.358 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.182 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M5 ;
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11] 
    ANTENNAPARTIALMETALAREA 0.023 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1012 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M4 ;
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10] 
    ANTENNAPARTIALMETALAREA 0.0615 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2706 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.1872 LAYER M4 ;
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.328 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.478 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1472 LAYER M4 ;
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2882 LAYER M2 ;
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 12.496 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 55.0704 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 2.646 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6864 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 247.854 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 1094.16 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.77994 LAYER VIA7 ;
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9152 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.386 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1424 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.858 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 47.8192 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 1.866 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2544 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 207.646 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 916.806 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA7 ;
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4768 LAYER M3 ;
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.222 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 31.8208 LAYER M6 ;
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3] 
    ANTENNAPARTIALMETALAREA 0.019 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0836 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0608 LAYER M3 ;
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2] 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.498 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2352 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.838 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 16.9312 LAYER M6 ;
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1] 
    ANTENNAPARTIALMETALAREA 0.051 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2244 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.706 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5504 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.378 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.3072 LAYER M4 ;
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0] 
    ANTENNAPARTIALMETALAREA 0.0225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.398 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1952 LAYER M3 ;
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.066 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M2 ;
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12] 
    ANTENNAPARTIALMETALAREA 0.0225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M3 ;
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.538 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8112 LAYER M4 ;
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.162 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M5 ;
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.006 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.2704 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.338 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9312 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.214 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0736 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M5 ; 
    ANTENNAMAXAREACAR 109.901 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 487.383 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA5 ;
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0285 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1694 LAYER M2 ;
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3568 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.996 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.8704 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 62.6675 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 279.557 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.666667 LAYER VIA4 ;
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.802 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.966 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2944 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.098 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.0752 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 193.768 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 855.663 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.33333 LAYER VIA6 ;
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.646 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6864 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.858 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 43.4192 LAYER M6 ;
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4] 
    ANTENNAPARTIALMETALAREA 1.0645 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6838 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.408 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M3 ;
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.506 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.178 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.4272 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 182.628 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 807.815 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA6 ;
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.422 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.222 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4208 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.638 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 42.4512 LAYER M6 ;
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.126 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.7984 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.318 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4432 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.198 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.5152 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 283.421 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1250.18 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6 ;
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0] 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.998 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.2352 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.34 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.584 LAYER M6 ;
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.171 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7524 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1395 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6578 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.166 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1744 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0471 LAYER M4 ; 
    ANTENNAMAXAREACAR 64.1062 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 284.153 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.06157 LAYER VIA4 ;
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4] 
    ANTENNAPARTIALMETALAREA 1.371 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.528 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.682 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0448 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 28.298 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 124.555 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.662 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 38.1568 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 LAYER M6 ; 
    ANTENNAMAXAREACAR 1681.52 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 7407.44 LAYER M6 ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VIA6 ;
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.9765 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2966 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.3342 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 104.29 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.504 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2616 LAYER M2 ;
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.811 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.759 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3836 LAYER M2 ;
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.2945 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3398 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6672 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0471 LAYER M4 ; 
    ANTENNAMAXAREACAR 65.1752 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 288.862 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.27389 LAYER VIA4 ;
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4] 
    ANTENNAPARTIALMETALAREA 1.09 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.84 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 17.8463 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 77.2958 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.138 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M3 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.8377 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 86.6926 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.1695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7458 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.638 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6512 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 65.65 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 290.51 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA4 ;
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.295 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.298 LAYER M2 ;
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.071 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3124 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.518 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7232 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 51.2844 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 227.832 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.809061 LAYER VIA4 ;
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0] 
    ANTENNAPARTIALMETALAREA 0.126 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5544 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.618 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.858 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6192 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 62.8378 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 277.955 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.402 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M5 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 69.3426 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 307.288 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA5 ;
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[15] 
    ANTENNAPARTIALMETALAREA 0.171 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7524 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9152 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.986 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.5824 LAYER M5 ;
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14] 
    ANTENNAPARTIALMETALAREA 0.111 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4884 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.338 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M4 ;
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13] 
    ANTENNAPARTIALMETALAREA 0.3455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5202 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.5888 LAYER M3 ;
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12] 
    ANTENNAPARTIALMETALAREA 0.097 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4268 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.618 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 4.982 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.9648 LAYER M5 ;
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11] 
    ANTENNAPARTIALMETALAREA 0.1115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4906 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.446 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0064 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 4.898 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5952 LAYER M5 ;
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10] 
    ANTENNAPARTIALMETALAREA 0.549 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4156 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0208 LAYER M3 ;
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4586 LAYER M2 ;
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8] 
    ANTENNAPARTIALMETALAREA 0.171 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7524 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 4.602 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.2928 LAYER M5 ;
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7] 
    ANTENNAPARTIALMETALAREA 0.4125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.815 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.738 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.0912 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 30.182 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 132.845 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.102 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 2.822 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 12.4608 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 413.421 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 1824.32 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.77994 LAYER VIA7 ;
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.467 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0548 LAYER M2 ;
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2945 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3398 LAYER M2 ;
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.686 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0624 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 14.4174 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 65.1486 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4 ;
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3] 
    ANTENNAPARTIALMETALAREA 0.741 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3044 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 11.3149 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 50.228 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.0379 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 67.2439 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.697 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 15.882 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 70.3232 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.1443 LAYER VIA2 ;
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1] 
    ANTENNAPARTIALMETALAREA 0.591 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6004 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.676 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0184 LAYER M2 ;
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13] 
    ANTENNAPARTIALMETALAREA 0.143 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6292 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.586 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.498 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6352 LAYER M4 ;
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12] 
    ANTENNAPARTIALMETALAREA 0.0745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3278 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.842 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6752 LAYER M4 ;
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.882 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9248 LAYER M3 ;
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.7445 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.9198 LAYER M2 ;
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9] 
    ANTENNAPARTIALMETALAREA 0.07 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.308 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M3 ;
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8] 
    ANTENNAPARTIALMETALAREA 1.1305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.566 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5344 LAYER M3 ;
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7] 
    ANTENNAPARTIALMETALAREA 0.23 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.012 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.986 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3824 LAYER M3 ;
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0265 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1606 LAYER M2 ;
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7808 LAYER M3 ;
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0226 LAYER M2 ;
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.426 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9184 LAYER M3 ;
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0394 LAYER M2 ;
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.063 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3212 LAYER M2 ;
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4158 LAYER M2 ;
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5015 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2506 LAYER M2 ;
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 1.05 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.62 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.392 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.2128 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.958 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 24.082 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 106.005 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.394 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 37.0656 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 385.62 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1701.7 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA6 ;
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7065 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1526 LAYER M2 ;
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.181 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2404 LAYER M2 ;
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.2955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7442 LAYER M2 ;
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.166 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7304 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.718 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.026 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5584 LAYER M4 ;
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.2975 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.353 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 77.1982 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 329.12 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA3 ;
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.357 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5708 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.942 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1888 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 91.8855 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 403.563 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA4 ;
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.2085 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9174 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.914 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.2512 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 199.654 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA3 ;
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 1.428 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2832 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.288 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.4947 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 206.757 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1] 
    ANTENNAPARTIALMETALAREA 1.1775 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.181 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.6272 LAYER M3 ;
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.571 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5124 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0608 LAYER M3 ;
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.6285 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7654 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.698 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1152 LAYER M3 ;
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.111 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4884 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.662 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9568 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.878 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7072 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 93.7443 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 414.893 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA5 ;
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.1185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.942 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.8768 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 85.2977 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 378.44 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.809061 LAYER VIA4 ;
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.713 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1812 LAYER M2 ;
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1] 
    ANTENNAPARTIALMETALAREA 2.9075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.793 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 138.67 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 612.79 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3 ;
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.351 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.23 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.856 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 77.8932 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 343.948 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.618 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1632 LAYER M4 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 130.256 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 575.767 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA4 ;
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5] 
    ANTENNAPARTIALMETALAREA 1.2255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3922 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.6352 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 126.975 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.471698 LAYER VIA3 ;
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4] 
    ANTENNAPARTIALMETALAREA 1.016 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4704 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.208 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.6032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.8307 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 224.081 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.209644 LAYER VIA3 ;
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3] 
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.406 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2304 LAYER M4 ;
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.391 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7204 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.176 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2184 LAYER M3 ;
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.7945 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4958 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.946 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 80.4215 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 353.042 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA3 ;
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.311 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2 ;
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13] 
    ANTENNAPARTIALMETALAREA 4.915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.67 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.406 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M3 ;
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12] 
    ANTENNAPARTIALMETALAREA 0.0315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1386 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.018 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5232 LAYER M4 ;
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.6785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8294 LAYER M2 ;
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.718 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M4 ;
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M3 ;
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.458 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.358 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M4 ;
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.3015 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.3266 LAYER M2 ;
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.246 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5264 LAYER M3 ;
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0604 LAYER M2 ;
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.758 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3792 LAYER M3 ;
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8048 LAYER M3 ;
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.418 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M4 ;
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done 
    ANTENNAPARTIALMETALAREA 0.226 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9944 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.6272 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 8.798 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 38.7552 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 3.386 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 14.9424 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M7 ; 
    ANTENNAMAXAREACAR 194.869 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 864.257 LAYER M7 ;
    ANTENNAMAXCUTCAR 2.77078 LAYER VIA7 ;
  END dsadc_conv_done
  PIN dsadc_en 
    ANTENNAPARTIALMETALAREA 0.272 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.258 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.1792 LAYER M5 ;
  END dsadc_en
  PIN dsadc_clk 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 17.864 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8264 LAYER M3 ;
  END dsadc_clk
  PIN dsadc_switch[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1318 LAYER M2 ;
  END dsadc_switch[2]
  PIN dsadc_switch[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.285 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.298 LAYER M2 ;
  END dsadc_switch[1]
  PIN dsadc_switch[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.155 LAYER M2 ;
  END dsadc_switch[0]
  PIN dac_en_pot 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0814 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.718 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.018 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1232 LAYER M5 ;
  END dac_en_pot
  PIN adc_ext_in 
    ANTENNAPARTIALMETALAREA 0.487 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1428 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.6608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.278 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6672 LAYER M5 ;
  END adc_ext_in
  PIN atp_en 
    ANTENNAPARTIALMETALAREA 0.9205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0502 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.6848 LAYER M3 ;
  END atp_en
  PIN atp_sel 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.377 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7028 LAYER M2 ;
  END atp_sel
  PIN adc_sel 
    ANTENNAPARTIALMETALAREA 0.1135 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4994 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.624 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0336 LAYER M5 ;
  END adc_sel
  PIN saradc_clk 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 66.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.4602 LAYER M3 ;
  END saradc_clk
  PIN saradc_rdy 
    ANTENNAPARTIALMETALAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.866 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8544 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M4 ; 
    ANTENNAMAXAREACAR 412.694 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1817.45 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.21402 LAYER VIA4 ;
  END saradc_rdy
  PIN saradc_rst 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.331 LAYER M2 ;
  END saradc_rst
  PIN saradc_data[9] 
    ANTENNAPARTIALMETALAREA 0.616 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7984 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 24.345 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 108.908 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2 ;
  END saradc_data[9]
  PIN saradc_data[8] 
    ANTENNAPARTIALMETALAREA 0.1515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3232 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M4 ; 
    ANTENNAMAXAREACAR 350.923 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1541.67 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.21402 LAYER VIA4 ;
  END saradc_data[8]
  PIN saradc_data[7] 
    ANTENNAPARTIALMETALAREA 0.4515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9866 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 6.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.5968 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 269.594 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1176.09 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[7]
  PIN saradc_data[6] 
    ANTENNAPARTIALMETALAREA 0.5065 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 7.678 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.8272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 315.661 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1367.38 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[6]
  PIN saradc_data[5] 
    ANTENNAPARTIALMETALAREA 0.5915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6026 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M4 ; 
    ANTENNAMAXAREACAR 407.085 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1791.7 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.21402 LAYER VIA4 ;
  END saradc_data[5]
  PIN saradc_data[4] 
    ANTENNAPARTIALMETALAREA 0.227 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9988 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.8575 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 52.217 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 469.886 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2045.97 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[4]
  PIN saradc_data[3] 
    ANTENNAPARTIALMETALAREA 0.3115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3706 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.418 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.8832 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 162.45 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 714.83 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END saradc_data[3]
  PIN saradc_data[2] 
    ANTENNAPARTIALMETALAREA 0.4065 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7886 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.6928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 404.502 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1777.65 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[2]
  PIN saradc_data[1] 
    ANTENNAPARTIALMETALAREA 1.1615 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1546 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.2608 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 400 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1759.7 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[1]
  PIN saradc_data[0] 
    ANTENNAPARTIALMETALAREA 0.3035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 7.498 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.0352 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 304.059 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1330.13 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END saradc_data[0]
END MCU

END LIBRARY
