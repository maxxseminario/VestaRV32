

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO MCU 
  PIN resetn_in 
    ANTENNAPARTIALMETALAREA 0.9625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.235 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.658 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9392 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 24.822 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 109.261 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 939.327 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4139.7 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6 ;
  END resetn_in
  PIN resetn_out 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.474 LAYER M2 ;
  END resetn_out
  PIN resetn_dir 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6365 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8446 LAYER M2 ;
  END resetn_dir
  PIN resetn_ren 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6378 LAYER M2 ;
  END resetn_ren
  PIN prt1_in[7] 
    ANTENNAPARTIALMETALAREA 0.1125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.495 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 607.666 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2675.52 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3 ;
  END prt1_in[7]
  PIN prt1_in[6] 
    ANTENNAPARTIALMETALAREA 21.6165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 95.1126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.3088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 112.847 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 494.349 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.734684 LAYER VIA3 ;
  END prt1_in[6]
  PIN prt1_in[5] 
    ANTENNAPARTIALMETALAREA 1.1725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.159 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.756 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.9024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1305 LAYER M3 ; 
    ANTENNAMAXAREACAR 102.335 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 450.859 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.93942 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 3.698 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3152 LAYER M4 ;
    ANTENNAGATEAREA 0.1941 LAYER M4 ; 
    ANTENNAMAXAREACAR 121.387 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 534.914 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.943396 LAYER VIA4 ;
  END prt1_in[5]
  PIN prt1_in[4] 
    ANTENNAPARTIALMETALAREA 0.0325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.143 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.66 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1305 LAYER M4 ; 
    ANTENNAMAXAREACAR 174.297 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 768.726 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 1.24593 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.466 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.6944 LAYER M5 ;
    ANTENNAGATEAREA 0.2577 LAYER M5 ; 
    ANTENNAMAXAREACAR 191.627 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 845.15 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.24593 LAYER VIA5 ;
  END prt1_in[4]
  PIN prt1_in[3] 
    ANTENNAPARTIALMETALAREA 0.176 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1936 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7622 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.64 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M4 ; 
    ANTENNAMAXAREACAR 18.0514 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 23.5577 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 0.419287 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 9.92 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.088 LAYER M5 ;
    ANTENNAGATEAREA 0.2544 LAYER M5 ; 
    ANTENNAMAXAREACAR 57.0451 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 75.9623 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.25786 LAYER VIA5 ;
  END prt1_in[3]
  PIN prt1_in[2] 
    ANTENNAPARTIALMETALAREA 4.6775 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.625 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.41 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0671 LAYER M3 ; 
    ANTENNAMAXAREACAR 172.381 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 758.73 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.894188 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.098 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8752 LAYER M4 ;
    ANTENNAGATEAREA 0.1709 LAYER M4 ; 
    ANTENNAMAXAREACAR 178.806 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 787.257 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.27669 LAYER VIA4 ;
  END prt1_in[2]
  PIN prt1_in[1] 
    ANTENNAPARTIALMETALAREA 13.3775 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.905 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.4928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.0464 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 264.02 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[1]
  PIN prt1_in[0] 
    ANTENNAPARTIALMETALAREA 24.0995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 106.038 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.1088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 LAYER M3 ; 
    ANTENNAMAXAREACAR 88.9885 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 392.049 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.542005 LAYER VIA3 ;
  END prt1_in[0]
  PIN prt1_out[7] 
    ANTENNAPARTIALMETALAREA 1.872 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2368 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.224 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.6736 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 33.562 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 147.717 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2242 LAYER M6 ; 
    ANTENNAMAXAREACAR 167.101 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 734.874 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.02592 LAYER VIA6 ;
  END prt1_out[7]
  PIN prt1_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.657 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 55.8228 LAYER M2 ;
  END prt1_out[6]
  PIN prt1_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.821 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
  END prt1_out[5]
  PIN prt1_out[4] 
    ANTENNAPARTIALMETALAREA 1.754 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7616 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.8048 LAYER M3 ;
  END prt1_out[4]
  PIN prt1_out[3] 
    ANTENNAPARTIALMETALAREA 0.956 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2064 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.4448 LAYER M3 ;
  END prt1_out[3]
  PIN prt1_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[2]
  PIN prt1_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[1]
  PIN prt1_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 52.426 LAYER M2 ;
  END prt1_out[0]
  PIN prt1_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.6015 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.2906 LAYER M2 ;
  END prt1_dir[7]
  PIN prt1_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.8415 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 52.1466 LAYER M2 ;
  END prt1_dir[6]
  PIN prt1_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.2035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.1834 LAYER M2 ;
  END prt1_dir[5]
  PIN prt1_dir[4] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[4]
  PIN prt1_dir[3] 
    ANTENNAPARTIALMETALAREA 0.6965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0646 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.022 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.9408 LAYER M3 ;
  END prt1_dir[3]
  PIN prt1_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
  END prt1_dir[2]
  PIN prt1_dir[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[1]
  PIN prt1_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.7745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.2958 LAYER M2 ;
  END prt1_dir[0]
  PIN prt1_ren[7] 
    ANTENNAPARTIALMETALAREA 0.1005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4422 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.486 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5824 LAYER M3 ;
  END prt1_ren[7]
  PIN prt1_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.3835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.9754 LAYER M2 ;
  END prt1_ren[6]
  PIN prt1_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.8275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 60.929 LAYER M2 ;
  END prt1_ren[5]
  PIN prt1_ren[4] 
    ANTENNAPARTIALMETALAREA 2.2785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0694 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.066 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.1344 LAYER M3 ;
  END prt1_ren[4]
  PIN prt1_ren[3] 
    ANTENNAPARTIALMETALAREA 0.5205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.618 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.3632 LAYER M3 ;
  END prt1_ren[3]
  PIN prt1_ren[2] 
    ANTENNAPARTIALMETALAREA 1.5455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.152 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.3568 LAYER M3 ;
  END prt1_ren[2]
  PIN prt1_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.3705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 54.5182 LAYER M2 ;
  END prt1_ren[1]
  PIN prt1_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.7305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.1022 LAYER M2 ;
  END prt1_ren[0]
  PIN prt2_in[7] 
    ANTENNAPARTIALMETALAREA 0.7735 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4474 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 8.45283 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 36.1022 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2 ;
  END prt2_in[7]
  PIN prt2_in[6] 
    ANTENNAPARTIALMETALAREA 0.7585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4254 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 23.0778 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 103.02 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.288184 LAYER VIA2 ;
  END prt2_in[6]
  PIN prt2_in[5] 
    ANTENNAPARTIALMETALAREA 0.9355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1162 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.426 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.6639 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 158.244 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.37037 LAYER VIA3 ;
  END prt2_in[5]
  PIN prt2_in[4] 
    ANTENNAPARTIALMETALAREA 0.8445 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7598 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 7.2728 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 31.6242 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2 ;
  END prt2_in[4]
  PIN prt2_in[3] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3916 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.64 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.08 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3816 LAYER M4 ; 
    ANTENNAMAXAREACAR 9.3864 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 12.586 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA4 ;
  END prt2_in[3]
  PIN prt2_in[2] 
    ANTENNAPARTIALMETALAREA 0.3155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.2448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 601.024 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2646.3 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3 ;
  END prt2_in[2]
  PIN prt2_in[1] 
    ANTENNAPARTIALMETALAREA 0.6755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9722 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2214 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.88347 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 16.4734 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0903342 LAYER VIA2 ;
  END prt2_in[1]
  PIN prt2_in[0] 
    ANTENNAPARTIALMETALAREA 0.3535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5994 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 4.72642 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 19.8758 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2 ;
  END prt2_in[0]
  PIN prt2_out[7] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.463 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0372 LAYER M2 ;
  END prt2_out[7]
  PIN prt2_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.701 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1284 LAYER M2 ;
  END prt2_out[6]
  PIN prt2_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.579 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6356 LAYER M2 ;
  END prt2_out[5]
  PIN prt2_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.717 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1988 LAYER M2 ;
  END prt2_out[4]
  PIN prt2_out[3] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2 ;
  END prt2_out[3]
  PIN prt2_out[2] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.408 LAYER M2 ;
  END prt2_out[2]
  PIN prt2_out[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.279 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2276 LAYER M2 ;
  END prt2_out[1]
  PIN prt2_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.292 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M2 ;
  END prt2_out[0]
  PIN prt2_dir[7] 
    ANTENNAPARTIALMETALAREA 0.4965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1846 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.026 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1584 LAYER M3 ;
  END prt2_dir[7]
  PIN prt2_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1086 LAYER M2 ;
  END prt2_dir[6]
  PIN prt2_dir[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1198 LAYER M2 ;
  END prt2_dir[5]
  PIN prt2_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3486 LAYER M2 ;
  END prt2_dir[4]
  PIN prt2_dir[3] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.642 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.0688 LAYER M3 ;
  END prt2_dir[3]
  PIN prt2_dir[2] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5365 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3606 LAYER M2 ;
  END prt2_dir[2]
  PIN prt2_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2 ;
  END prt2_dir[1]
  PIN prt2_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3166 LAYER M2 ;
  END prt2_dir[0]
  PIN prt2_ren[7] 
    ANTENNAPARTIALMETALAREA 0.7035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.042 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.8288 LAYER M3 ;
  END prt2_ren[7]
  PIN prt2_ren[6] 
    ANTENNAPARTIALMETALAREA 0.447 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9668 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.5895 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6378 LAYER M3 ;
  END prt2_ren[6]
  PIN prt2_ren[5] 
    ANTENNAPARTIALMETALAREA 0.6105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6862 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.946 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.0064 LAYER M3 ;
  END prt2_ren[5]
  PIN prt2_ren[4] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3034 LAYER M2 ;
  END prt2_ren[4]
  PIN prt2_ren[3] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.362 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M4 ;
  END prt2_ren[3]
  PIN prt2_ren[2] 
    ANTENNAPARTIALMETALAREA 0.667 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9348 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.4095 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.6458 LAYER M3 ;
  END prt2_ren[2]
  PIN prt2_ren[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3295 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4938 LAYER M2 ;
  END prt2_ren[1]
  PIN prt2_ren[0] 
    ANTENNAPARTIALMETALAREA 0.6275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.761 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.126 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3984 LAYER M3 ;
  END prt2_ren[0]
  PIN prt3_in[7] 
    ANTENNAPARTIALMETALAREA 18.6195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 82.0138 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 690.83 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3040.15 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.738007 LAYER VIA2 ;
  END prt3_in[7]
  PIN prt3_in[6] 
    ANTENNAPARTIALMETALAREA 15.5145 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 68.3078 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.318 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.6432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 527.764 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2299.04 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[6]
  PIN prt3_in[5] 
    ANTENNAPARTIALMETALAREA 7.2565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.9286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.678 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.2272 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.814 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0256 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 28.4786 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 127.654 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA4 ;
  END prt3_in[5]
  PIN prt3_in[4] 
    ANTENNAPARTIALMETALAREA 0.2925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.287 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.042 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.2288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.382 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.3248 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M5 ; 
    ANTENNAMAXAREACAR 50.1752 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 221.435 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.876988 LAYER VIA5 ;
  END prt3_in[4]
  PIN prt3_in[3] 
    ANTENNAPARTIALMETALAREA 0.1755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7722 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 17.754 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.2496 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 LAYER M3 ; 
    ANTENNAMAXAREACAR 149.102 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 657.553 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA3 ;
  END prt3_in[3]
  PIN prt3_in[2] 
    ANTENNAPARTIALMETALAREA 2.1515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.5546 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 419.105 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1847.48 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3 ;
  END prt3_in[2]
  PIN prt3_in[1] 
    ANTENNAPARTIALMETALAREA 23.4935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 103.415 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.1488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 193.225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 828.399 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[1]
  PIN prt3_in[0] 
    ANTENNAPARTIALMETALAREA 0.0355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1562 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 300.444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1307.52 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt3_in[0]
  PIN prt3_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.821 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.3444 LAYER M2 ;
  END prt3_out[7]
  PIN prt3_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.394 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.1776 LAYER M2 ;
  END prt3_out[6]
  PIN prt3_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.137 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6468 LAYER M2 ;
  END prt3_out[5]
  PIN prt3_out[4] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.085 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.418 LAYER M2 ;
  END prt3_out[4]
  PIN prt3_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3124 LAYER M2 ;
  END prt3_out[3]
  PIN prt3_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.456 LAYER M2 ;
  END prt3_out[2]
  PIN prt3_out[1] 
    ANTENNAPARTIALMETALAREA 1.392 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1248 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.246 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5264 LAYER M3 ;
  END prt3_out[1]
  PIN prt3_out[0] 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.664 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.082 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8048 LAYER M4 ;
  END prt3_out[0]
  PIN prt3_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.1775 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 62.513 LAYER M2 ;
  END prt3_dir[7]
  PIN prt3_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 7.4595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.9098 LAYER M2 ;
  END prt3_dir[6]
  PIN prt3_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt3_dir[5]
  PIN prt3_dir[4] 
    ANTENNAPARTIALMETALAREA 0.3965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7446 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.0928 LAYER M3 ;
  END prt3_dir[4]
  PIN prt3_dir[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt3_dir[3]
  PIN prt3_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.1165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6446 LAYER M2 ;
  END prt3_dir[2]
  PIN prt3_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.8745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.1358 LAYER M2 ;
  END prt3_dir[1]
  PIN prt3_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.9255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0042 LAYER M2 ;
  END prt3_dir[0]
  PIN prt3_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.3655 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.9402 LAYER M2 ;
  END prt3_ren[7]
  PIN prt3_ren[6] 
    ANTENNAPARTIALMETALAREA 4.7425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.911 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.926 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9184 LAYER M3 ;
  END prt3_ren[6]
  PIN prt3_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.3415 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0346 LAYER M2 ;
  END prt3_ren[5]
  PIN prt3_ren[4] 
    ANTENNAPARTIALMETALAREA 0.4405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9382 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.6992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0582 LAYER M3 ; 
    ANTENNAMAXAREACAR 199.73 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 879.533 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.515464 LAYER VIA3 ;
  END prt3_ren[4]
  PIN prt3_ren[3] 
    ANTENNAPARTIALMETALAREA 0.4075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.793 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.984 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.0176 LAYER M3 ;
  END prt3_ren[3]
  PIN prt3_ren[2] 
    ANTENNAPARTIALMETALAREA 6.4255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.3162 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.882 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9248 LAYER M3 ;
  END prt3_ren[2]
  PIN prt3_ren[1] 
    ANTENNAPARTIALMETALAREA 11.2805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.6342 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.1568 LAYER M3 ;
  END prt3_ren[1]
  PIN prt3_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.6835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8954 LAYER M2 ;
  END prt3_ren[0]
  PIN prt4_in[7] 
    ANTENNAPARTIALMETALAREA 1.5555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 25.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 112.27 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 952.472 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4189.52 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt4_in[7]
  PIN prt4_in[6] 
    ANTENNAPARTIALMETALAREA 0.5355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3562 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 18.518 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 81.5232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 687.946 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3028.49 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3 ;
  END prt4_in[6]
  PIN prt4_in[5] 
    ANTENNAPARTIALMETALAREA 1.2385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4494 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.664 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.0096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M3 ; 
    ANTENNAMAXAREACAR 303.687 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1325.86 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.618 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M4 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 309.641 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1352.48 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA4 ;
  END prt4_in[5]
  PIN prt4_in[4] 
    ANTENNAPARTIALMETALAREA 7.0185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.8814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.498 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6352 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 7.738 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.0912 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M7 ; 
    ANTENNAMAXAREACAR 68.5396 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 304.614 LAYER M7 ;
    ANTENNAMAXCUTCAR 2.74606 LAYER VIA7 ;
  END prt4_in[4]
  PIN prt4_in[3] 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 16.826 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 74.0784 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M6 ; 
    ANTENNAMAXAREACAR 203.959 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 898.844 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.66205 LAYER VIA6 ;
  END prt4_in[3]
  PIN prt4_in[2] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 7.442 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.7888 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 16.286 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 71.7024 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M6 ; 
    ANTENNAMAXAREACAR 215.347 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 948.455 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.39104 LAYER VIA6 ;
  END prt4_in[2]
  PIN prt4_in[1] 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 648.28 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2845.08 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.69004 LAYER VIA6 ;
  END prt4_in[1]
  PIN prt4_in[0] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8528 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 15.822 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 69.6608 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 624.133 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2746.24 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.69004 LAYER VIA6 ;
  END prt4_in[0]
  PIN prt4_out[7] 
    ANTENNAPARTIALMETALAREA 5.292 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8806 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 82.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.08 LAYER M3 ;
  END prt4_out[7]
  PIN prt4_out[6] 
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 44.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.7542 LAYER M3 ;
  END prt4_out[6]
  PIN prt4_out[5] 
    ANTENNAPARTIALMETALAREA 0.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5654 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.592 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.2272 LAYER M3 ;
  END prt4_out[5]
  PIN prt4_out[4] 
    ANTENNAPARTIALMETALAREA 0.446 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4906 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.808 LAYER M3 ;
  END prt4_out[4]
  PIN prt4_out[3] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.0448 LAYER M3 ;
  END prt4_out[3]
  PIN prt4_out[2] 
    ANTENNAPARTIALMETALAREA 0.499 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1956 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.6384 LAYER M3 ;
  END prt4_out[2]
  PIN prt4_out[1] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.962 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 74.6768 LAYER M6 ;
  END prt4_out[1]
  PIN prt4_out[0] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[0]
  PIN prt4_dir[7] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1946 LAYER M2 ;
  END prt4_dir[7]
  PIN prt4_dir[6] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1946 LAYER M2 ;
  END prt4_dir[6]
  PIN prt4_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7358 LAYER M2 ;
  END prt4_dir[5]
  PIN prt4_dir[4] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2782 LAYER M2 ;
  END prt4_dir[4]
  PIN prt4_dir[3] 
    ANTENNAPARTIALMETALAREA 0.6965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0646 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.546 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0464 LAYER M3 ;
  END prt4_dir[3]
  PIN prt4_dir[2] 
    ANTENNAPARTIALMETALAREA 0.3565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5686 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.2384 LAYER M3 ;
  END prt4_dir[2]
  PIN prt4_dir[1] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 17.122 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 75.3808 LAYER M6 ;
  END prt4_dir[1]
  PIN prt4_dir[0] 
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6 ;
  END prt4_dir[0]
  PIN prt4_ren[7] 
    ANTENNAPARTIALMETALAREA 1.207 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3108 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.5255 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.1562 LAYER M3 ;
  END prt4_ren[7]
  PIN prt4_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.9475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.257 LAYER M2 ;
  END prt4_ren[6]
  PIN prt4_ren[5] 
    ANTENNAPARTIALMETALAREA 0.7105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1262 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.626 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.5984 LAYER M3 ;
  END prt4_ren[5]
  PIN prt4_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.4035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.8634 LAYER M2 ;
  END prt4_ren[4]
  PIN prt4_ren[3] 
    ANTENNAPARTIALMETALAREA 0.9235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0634 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.318 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0432 LAYER M3 ;
  END prt4_ren[3]
  PIN prt4_ren[2] 
    ANTENNAPARTIALMETALAREA 0.2805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2342 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.246 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.3264 LAYER M3 ;
  END prt4_ren[2]
  PIN prt4_ren[1] 
    ANTENNAPARTIALMETALAREA 0.8035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.366 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 72.0544 LAYER M6 ;
  END prt4_ren[1]
  PIN prt4_ren[0] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 17.142 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 75.4688 LAYER M6 ;
  END prt4_ren[0]
  PIN use_dac_glb_bias 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2022 LAYER M2 ;
  END use_dac_glb_bias
  PIN en_bias_buf 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.377 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7028 LAYER M2 ;
  END en_bias_buf
  PIN en_bias_gen 
    ANTENNAPARTIALMETALAREA 0.261 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1484 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.422 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10.598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 46.6752 LAYER M4 ;
  END en_bias_gen
  PIN BIAS_ADJ[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.354 LAYER M2 ;
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.318 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4432 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.022 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3408 LAYER M6 ;
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.3065 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8366 LAYER M2 ;
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.378 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7072 LAYER M3 ;
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0645 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3278 LAYER M2 ;
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.558 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.758 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1792 LAYER M4 ;
  END BIAS_DBP[13]
  PIN BIAS_DBP[12] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.702 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.798 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3552 LAYER M4 ;
  END BIAS_DBP[12]
  PIN BIAS_DBP[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DBP[11]
  PIN BIAS_DBP[10] 
    ANTENNAPARTIALMETALAREA 0.0705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3102 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.606 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1104 LAYER M3 ;
  END BIAS_DBP[10]
  PIN BIAS_DBP[9] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M3 ;
  END BIAS_DBP[9]
  PIN BIAS_DBP[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9558 LAYER M2 ;
  END BIAS_DBP[8]
  PIN BIAS_DBP[7] 
    ANTENNAPARTIALMETALAREA 0.487 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1428 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.942 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1888 LAYER M3 ;
  END BIAS_DBP[7]
  PIN BIAS_DBP[6] 
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.398 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1952 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.218 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.0032 LAYER M6 ;
  END BIAS_DBP[6]
  PIN BIAS_DBP[5] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.598 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0752 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.038 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.8112 LAYER M4 ;
  END BIAS_DBP[5]
  PIN BIAS_DBP[4] 
    ANTENNAPARTIALMETALAREA 0.2635 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1594 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9168 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.378 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1072 LAYER M4 ;
  END BIAS_DBP[4]
  PIN BIAS_DBP[3] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.666 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3744 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.878 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.3072 LAYER M4 ;
  END BIAS_DBP[3]
  PIN BIAS_DBP[2] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.418 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2832 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.758 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 51.7792 LAYER M6 ;
  END BIAS_DBP[2]
  PIN BIAS_DBP[1] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9872 LAYER M3 ;
  END BIAS_DBP[1]
  PIN BIAS_DBP[0] 
    ANTENNAPARTIALMETALAREA 0.1845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8558 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M3 ;
  END BIAS_DBP[0]
  PIN BIAS_DBN[13] 
    ANTENNAPARTIALMETALAREA 7.666 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.7744 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.046 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6464 LAYER M3 ;
  END BIAS_DBN[13]
  PIN BIAS_DBN[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 7.1475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.493 LAYER M2 ;
  END BIAS_DBN[12]
  PIN BIAS_DBN[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 7.082 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.2928 LAYER M2 ;
  END BIAS_DBN[11]
  PIN BIAS_DBN[10] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0655 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3322 LAYER M2 ;
  END BIAS_DBN[10]
  PIN BIAS_DBN[9] 
    ANTENNAPARTIALMETALAREA 0.129 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5676 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
  END BIAS_DBN[9]
  PIN BIAS_DBN[8] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9392 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.968 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.658 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.1392 LAYER M4 ;
  END BIAS_DBN[8]
  PIN BIAS_DBN[7] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M4 ;
  END BIAS_DBN[7]
  PIN BIAS_DBN[6] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.398 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7952 LAYER M3 ;
  END BIAS_DBN[6]
  PIN BIAS_DBN[5] 
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 8.842 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.9488 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 1.222 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4208 LAYER M7 ;
  END BIAS_DBN[5]
  PIN BIAS_DBN[4] 
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.698 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5152 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.178 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4272 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 5.338 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.5312 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 2.686 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8624 LAYER M7 ;
  END BIAS_DBN[4]
  PIN BIAS_DBN[3] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.962 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2768 LAYER M3 ;
  END BIAS_DBN[3]
  PIN BIAS_DBN[2] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.218 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 36.2032 LAYER M6 ;
  END BIAS_DBN[2]
  PIN BIAS_DBN[1] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.996 LAYER M3 ;
  END BIAS_DBN[1]
  PIN BIAS_DBN[0] 
    ANTENNAPARTIALMETALAREA 0.4335 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9514 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2128 LAYER M3 ;
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13] 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.338 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.538 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4112 LAYER M4 ;
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2335 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0714 LAYER M2 ;
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.21 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.968 LAYER M2 ;
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10] 
    ANTENNAPARTIALMETALAREA 0.0615 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2706 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.098 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2752 LAYER M4 ;
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5232 LAYER M3 ;
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8] 
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4448 LAYER M3 ;
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7] 
    ANTENNAPARTIALMETALAREA 0.57 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1008 LAYER M3 ;
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M4 ;
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.277 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7068 LAYER M2 ;
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.258 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.282 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6848 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.218 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.0032 LAYER M6 ;
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.722 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.778 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.0672 LAYER M4 ;
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.3275 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.485 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.262 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3968 LAYER M4 ;
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.802 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.7728 LAYER M4 ;
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0] 
    ANTENNAPARTIALMETALAREA 0.1605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7502 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.0992 LAYER M4 ;
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.018 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5232 LAYER M3 ;
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12] 
    ANTENNAPARTIALMETALAREA 0.1085 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4774 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.982 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.1648 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.882 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 39.1248 LAYER M6 ;
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.398 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7952 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.106 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M5 ;
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10] 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.458 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 37.2592 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 213.761 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 943.53 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9] 
    ANTENNAPARTIALMETALAREA 0.101 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4884 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.638 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8512 LAYER M3 ;
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.546 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8464 LAYER M3 ;
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9152 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.782 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.2848 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.946 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 43.8064 LAYER M6 ;
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6175 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.761 LAYER M2 ;
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5] 
    ANTENNAPARTIALMETALAREA 0.064 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2816 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.086 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4224 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.958 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 39.4592 LAYER M6 ;
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4] 
    ANTENNAPARTIALMETALAREA 1.8595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2258 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.398 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 36.9952 LAYER M6 ;
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3] 
    ANTENNAPARTIALMETALAREA 0.474 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4784 LAYER M3 ;
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2] 
    ANTENNAPARTIALMETALAREA 0.0615 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2706 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1808 LAYER M3 ;
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1] 
    ANTENNAPARTIALMETALAREA 0.023 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1012 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.958 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M3 ;
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0] 
    ANTENNAPARTIALMETALAREA 0.0195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.458 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0592 LAYER M3 ;
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.333 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5092 LAYER M2 ;
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.639 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8996 LAYER M2 ;
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.256 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M2 ;
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.707 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1988 LAYER M2 ;
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.556 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.17 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 36.4087 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 161.911 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4 ;
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3046 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.19 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.324 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.798 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5552 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 24.4986 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 109.117 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA5 ;
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.095 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.806 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5904 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 42.9113 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 189.498 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA4 ;
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.6265 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7566 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.206 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.7504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.0167 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 176.99 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.806 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5904 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.442 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3888 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M5 ; 
    ANTENNAMAXAREACAR 29.59 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 126.83 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA5 ;
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1] 
    ANTENNAPARTIALMETALAREA 1.0335 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5474 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.51 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 44.6177 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 197.074 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0] 
    ANTENNAPARTIALMETALAREA 1.186 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.308 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.4163 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.554 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[16] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5804 LAYER M2 ;
  END BIAS_TIA_G_POT[16]
  PIN BIAS_TIA_G_POT[15] 
    ANTENNAPARTIALMETALAREA 0.1165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.962 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2768 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 8.74 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 38.544 LAYER M5 ;
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14] 
    ANTENNAPARTIALMETALAREA 0.051 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2244 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.622 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 24.7808 LAYER M5 ;
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13] 
    ANTENNAPARTIALMETALAREA 0.3085 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.818 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0432 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 4.338 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.1312 LAYER M5 ;
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12] 
    ANTENNAPARTIALMETALAREA 0.211 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9284 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.738 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6912 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 4.082 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.0048 LAYER M5 ;
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11] 
    ANTENNAPARTIALMETALAREA 0.5945 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6158 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.146 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4864 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.758 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7792 LAYER M5 ;
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10] 
    ANTENNAPARTIALMETALAREA 0.385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.694 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 6.422 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 28.3008 LAYER M5 ;
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9] 
    ANTENNAPARTIALMETALAREA 0.3235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4234 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.702 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1328 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.862 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 25.8368 LAYER M5 ;
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8] 
    ANTENNAPARTIALMETALAREA 0.211 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9284 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.878 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9072 LAYER M4 ;
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3442 LAYER M2 ;
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6] 
    ANTENNAPARTIALMETALAREA 0.547 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.836 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.5664 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 60.168 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 264.915 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 14.822 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 65.2608 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 257.541 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1130.52 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5] 
    ANTENNAPARTIALMETALAREA 0.1585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6974 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.142 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.75 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.144 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 41.8056 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 185.657 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA4 ;
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4] 
    ANTENNAPARTIALMETALAREA 3.0805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.5542 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 45.074 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 198.133 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.426 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9184 LAYER M3 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 51.2211 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 225.815 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3] 
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0945 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4598 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.942 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1888 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M5 ; 
    ANTENNAMAXAREACAR 19.6122 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 89.2756 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA5 ;
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2] 
    ANTENNAPARTIALMETALAREA 0.051 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2244 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.356 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.11 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 155.561 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1] 
    ANTENNAPARTIALMETALAREA 0.1915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8426 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.478 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1472 LAYER M3 ;
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0] 
    ANTENNAPARTIALMETALAREA 0.077 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3388 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1648 LAYER M3 ;
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.198 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9152 LAYER M3 ;
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12] 
    ANTENNAPARTIALMETALAREA 0.2345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0318 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3 ;
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11] 
    ANTENNAPARTIALMETALAREA 0.069 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.4595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5098 LAYER M2 ;
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.198 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3152 LAYER M4 ;
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8] 
    ANTENNAPARTIALMETALAREA 0.1925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.847 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.686 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0624 LAYER M3 ;
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7] 
    ANTENNAPARTIALMETALAREA 0.07 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.308 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.626 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7984 LAYER M3 ;
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6] 
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6608 LAYER M3 ;
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3 ;
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.692 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M2 ;
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2] 
    ANTENNAPARTIALMETALAREA 0.0285 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1254 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.119 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5676 LAYER M2 ;
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4158 LAYER M2 ;
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.022 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.9329 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 166.416 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.33 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.452 LAYER M2 ;
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.6445 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8358 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.002 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4528 LAYER M3 ;
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.851 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.938 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.3846 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 142.309 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1] 
    ANTENNAPARTIALMETALAREA 1.071 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7124 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.718 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2032 LAYER M3 ;
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.738 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2912 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1135 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9434 LAYER M2 ;
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.171 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7524 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.108 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5192 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.886 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9424 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 87.8649 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 378.828 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA4 ;
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3] 
    ANTENNAPARTIALMETALAREA 1.4735 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5274 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M2 ; 
    ANTENNAMAXAREACAR 39.8062 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 168.913 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.906 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0304 LAYER M3 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 54.4664 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 234.129 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA3 ;
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.934 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1536 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.738 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.3062 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 142.1 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.2065 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3526 LAYER M2 ;
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.517 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3188 LAYER M2 ;
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.027 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1188 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0705 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3542 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.958 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M5 ; 
    ANTENNAMAXAREACAR 73.3625 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 326.861 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.26537 LAYER VIA5 ;
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.667 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9348 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 69.9968 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 309.204 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3 ;
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.135 LAYER M2 ;
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.209 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9196 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.082 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8048 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 38.6958 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 171.968 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.809061 LAYER VIA4 ;
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1] 
    ANTENNAPARTIALMETALAREA 1.1465 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0446 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.778 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.8672 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.546 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4464 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 LAYER M4 ; 
    ANTENNAMAXAREACAR 18.2467 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 82.3111 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.11111 LAYER VIA4 ;
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.851 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.2201 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 183.074 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.478 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1472 LAYER M3 ;
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.779 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5156 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.766 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4144 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.202 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 23.538 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 103.611 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.166 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 1.522 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7408 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M7 ; 
    ANTENNAMAXAREACAR 166.311 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 733.676 LAYER M7 ;
    ANTENNAMAXCUTCAR 3.8835 LAYER VIA7 ;
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.726 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2384 LAYER M2 ;
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.129 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5676 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.382 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2304 LAYER M4 ; 
    ANTENNAMAXAREACAR 56.39 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 248.344 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.260417 LAYER VIA4 ;
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.6115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6906 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.586 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0224 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ; 
    ANTENNAMAXAREACAR 66.0894 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 288.938 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.33333 LAYER VIA3 ;
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0] 
    ANTENNAPARTIALMETALAREA 1.239 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4956 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.9729 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 157.531 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA3 ;
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.95 LAYER M2 ;
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12] 
    ANTENNAPARTIALMETALAREA 0.0315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1386 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1016 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.484 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.898 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9952 LAYER M4 ;
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11] 
    ANTENNAPARTIALMETALAREA 0.129 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5676 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.1205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6182 LAYER M2 ;
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.338 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3312 LAYER M4 ;
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6] 
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M3 ;
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.582 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6048 LAYER M3 ;
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.692 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.546 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4464 LAYER M3 ;
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3] 
    ANTENNAPARTIALMETALAREA 5.583 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.6092 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.192 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.1328 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 119.881 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 528.165 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.2886 LAYER VIA3 ;
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2] 
    ANTENNAPARTIALMETALAREA 0.2165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9526 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.866 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8544 LAYER M3 ;
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1] 
    ANTENNAPARTIALMETALAREA 0.071 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3124 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3088 LAYER M3 ;
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0875 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.429 LAYER M2 ;
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done 
    ANTENNAPARTIALMETALAREA 0.042 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1848 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.378 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.3072 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 3.646 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0864 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M7 ; 
    ANTENNAMAXAREACAR 181.385 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 800.035 LAYER M7 ;
    ANTENNAMAXCUTCAR 3.02267 LAYER VIA7 ;
  END dsadc_conv_done
  PIN dsadc_en 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.474 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1296 LAYER M2 ;
  END dsadc_en
  PIN dsadc_clk 
    ANTENNAPARTIALMETALAREA 1.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.984 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.6584 LAYER M3 ;
  END dsadc_clk
  PIN dsadc_switch[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.526 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M2 ;
  END dsadc_switch[2]
  PIN dsadc_switch[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.268 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M2 ;
  END dsadc_switch[1]
  PIN dsadc_switch[0] 
    ANTENNAPARTIALMETALAREA 0.3185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4014 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.406 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2304 LAYER M3 ;
  END dsadc_switch[0]
  PIN dac_en_pot 
    ANTENNAPARTIALMETALAREA 0.251 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1044 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.3185 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8454 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.298 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1552 LAYER M5 ;
  END dac_en_pot
  PIN adc_ext_in 
    ANTENNAPARTIALMETALAREA 1.453 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4372 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9968 LAYER M3 ;
  END adc_ext_in
  PIN atp_en 
    ANTENNAPARTIALMETALAREA 0.1645 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7238 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.038 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.0112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.238 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M4 ;
  END atp_en
  PIN atp_sel 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.377 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7028 LAYER M2 ;
  END atp_sel
  PIN adc_sel 
    ANTENNAPARTIALMETALAREA 0.1535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9944 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.398 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7952 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 2.922 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9008 LAYER M7 ;
  END adc_sel
  PIN saradc_clk 
    ANTENNAPARTIALMETALAREA 1.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 69.422 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.7162 LAYER M3 ;
  END saradc_clk
  PIN saradc_rdy 
    ANTENNAPARTIALMETALAREA 0.6425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.827 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0676 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.702 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5328 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.278 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6672 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.628 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8512 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 1.486 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5824 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M7 ; 
    ANTENNAMAXAREACAR 131.28 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 574.496 LAYER M7 ;
    ANTENNAMAXCUTCAR 3.45821 LAYER VIA7 ;
  END saradc_rdy
  PIN saradc_rst 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1726 LAYER M2 ;
  END saradc_rst
  PIN saradc_data[9] 
    ANTENNAPARTIALMETALAREA 0.3025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.331 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.778 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.0672 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.422 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.9008 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0269 LAYER M5 ; 
    ANTENNAMAXAREACAR 249.108 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1098.88 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.97398 LAYER VIA5 ;
  END saradc_data[9]
  PIN saradc_data[8] 
    ANTENNAPARTIALMETALAREA 0.6425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.827 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.826 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.8784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 240.73 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1057.08 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END saradc_data[8]
  PIN saradc_data[7] 
    ANTENNAPARTIALMETALAREA 0.7845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4958 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 7.022 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.9408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 199.068 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 872.861 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END saradc_data[7]
  PIN saradc_data[6] 
    ANTENNAPARTIALMETALAREA 0.567 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4948 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.2815 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.702 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 60.3328 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 611.267 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2678.84 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[6]
  PIN saradc_data[5] 
    ANTENNAPARTIALMETALAREA 0.9155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0282 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.7488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 236.549 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1038.5 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END saradc_data[5]
  PIN saradc_data[4] 
    ANTENNAPARTIALMETALAREA 0.651 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8644 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.2935 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.9354 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 9.478 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 41.7472 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 451.414 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1984.83 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.85714 LAYER VIA5 ;
  END saradc_data[4]
  PIN saradc_data[3] 
    ANTENNAPARTIALMETALAREA 0.8915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9226 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.958 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 12.116 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 53.3984 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 541.227 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2373.31 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[3]
  PIN saradc_data[2] 
    ANTENNAPARTIALMETALAREA 0.8425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.707 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.022 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.1408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 310 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1364.05 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END saradc_data[2]
  PIN saradc_data[1] 
    ANTENNAPARTIALMETALAREA 0.7225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.179 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.858 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8192 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 11.338 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 49.9312 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.546 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4464 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 1.622 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1808 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M7 ; 
    ANTENNAMAXAREACAR 126.369 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 549.731 LAYER M7 ;
    ANTENNAMAXCUTCAR 4.89796 LAYER VIA7 ;
  END saradc_data[1]
  PIN saradc_data[0] 
    ANTENNAPARTIALMETALAREA 0.2395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0538 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.0464 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 9.342 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 41.1488 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6 ; 
    ANTENNAMAXAREACAR 209.635 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 910.188 LAYER M6 ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6 ;
  END saradc_data[0]
END MCU

END LIBRARY
