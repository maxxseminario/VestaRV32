/home/mseminario2/chips/myshkin/ic/abstracts/myshkin_abs/OscillatorCurrentStarved/OscillatorCurrentStarved.lef