

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO MCU 
  PIN resetn_in 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 25.922 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 114.101 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 974.013 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4292.32 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6 ;
  END resetn_in
  PIN resetn_out 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.474 LAYER M2 ;
  END resetn_out
  PIN resetn_dir 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6654 LAYER M2 ;
  END resetn_dir
  PIN resetn_ren 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1086 LAYER M2 ;
  END resetn_ren
  PIN prt1_in[7] 
    ANTENNAPARTIALMETALAREA 0.1125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.495 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 583.026 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2565.02 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt1_in[7]
  PIN prt1_in[6] 
    ANTENNAPARTIALMETALAREA 14.1925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 62.447 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.658 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.9392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 235.808 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1018.15 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt1_in[6]
  PIN prt1_in[5] 
    ANTENNAPARTIALMETALAREA 7.0325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.943 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.526 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.5584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 173.829 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 748.569 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END prt1_in[5]
  PIN prt1_in[4] 
    ANTENNAPARTIALMETALAREA 7.0125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.855 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.684 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.2976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2577 LAYER M3 ; 
    ANTENNAMAXAREACAR 64.8822 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 284.876 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.935444 LAYER VIA3 ;
  END prt1_in[4]
  PIN prt1_in[3] 
    ANTENNAPARTIALMETALAREA 0.176 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1936 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.964 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2364 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 19.36 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.648 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER M5 ; 
    ANTENNAMAXAREACAR 146.799 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 177.903 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.88679 LAYER VIA5 ;
  END prt1_in[3]
  PIN prt1_in[2] 
    ANTENNAPARTIALMETALAREA 5.0155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.0682 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.178 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.2272 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.916 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5184 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1776 LAYER M4 ; 
    ANTENNAMAXAREACAR 63.2544 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 281.931 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.43902 LAYER VIA4 ;
  END prt1_in[2]
  PIN prt1_in[1] 
    ANTENNAPARTIALMETALAREA 1.2935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.092 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.6928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.9202 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 166.811 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[1]
  PIN prt1_in[0] 
    ANTENNAPARTIALMETALAREA 7.8195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.4058 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.5568 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 218.144 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 959.649 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[0]
  PIN prt1_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 8.214 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.1856 LAYER M2 ;
  END prt1_out[7]
  PIN prt1_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
  END prt1_out[6]
  PIN prt1_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.043 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.6772 LAYER M2 ;
  END prt1_out[5]
  PIN prt1_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[4]
  PIN prt1_out[3] 
    ANTENNAPARTIALMETALAREA 0.976 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2944 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.5088 LAYER M3 ;
  END prt1_out[3]
  PIN prt1_out[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[2]
  PIN prt1_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[1]
  PIN prt1_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 10.699 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 47.1636 LAYER M2 ;
  END prt1_out[0]
  PIN prt1_dir[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[7]
  PIN prt1_dir[6] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
  END prt1_dir[6]
  PIN prt1_dir[5] 
    ANTENNAPARTIALMETALAREA 5.2345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0758 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.9904 LAYER M3 ;
  END prt1_dir[5]
  PIN prt1_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
  END prt1_dir[4]
  PIN prt1_dir[3] 
    ANTENNAPARTIALMETALAREA 0.7365 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2406 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.006 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.8704 LAYER M3 ;
  END prt1_dir[3]
  PIN prt1_dir[2] 
    ANTENNAPARTIALMETALAREA 5.2155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.9482 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.898 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.1952 LAYER M3 ;
  END prt1_dir[2]
  PIN prt1_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3486 LAYER M2 ;
  END prt1_dir[1]
  PIN prt1_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.5345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.8398 LAYER M2 ;
  END prt1_dir[0]
  PIN prt1_ren[7] 
    ANTENNAPARTIALMETALAREA 0.9605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2262 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.426 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3184 LAYER M3 ;
  END prt1_ren[7]
  PIN prt1_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.4255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.2042 LAYER M2 ;
  END prt1_ren[6]
  PIN prt1_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2 ;
  END prt1_ren[5]
  PIN prt1_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5962 LAYER M2 ;
  END prt1_ren[4]
  PIN prt1_ren[3] 
    ANTENNAPARTIALMETALAREA 0.1205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5302 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.802 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1728 LAYER M3 ;
  END prt1_ren[3]
  PIN prt1_ren[2] 
    ANTENNAPARTIALMETALAREA 4.5655 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.1322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.5408 LAYER M3 ;
  END prt1_ren[2]
  PIN prt1_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.5305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.8222 LAYER M2 ;
  END prt1_ren[1]
  PIN prt1_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.5305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.8222 LAYER M2 ;
  END prt1_ren[0]
  PIN prt2_in[7] 
    ANTENNAPARTIALMETALAREA 0.7505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3462 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0671 LAYER M2 ; 
    ANTENNAMAXAREACAR 15.8756 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 68.1639 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.298063 LAYER VIA2 ;
  END prt2_in[7]
  PIN prt2_in[6] 
    ANTENNAPARTIALMETALAREA 0.5555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 18.9193 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 83.7118 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END prt2_in[6]
  PIN prt2_in[5] 
    ANTENNAPARTIALMETALAREA 0.731 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M3 ; 
    ANTENNAMAXAREACAR 130.435 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 562.465 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.63265 LAYER VIA3 ;
  END prt2_in[5]
  PIN prt2_in[4] 
    ANTENNAPARTIALMETALAREA 0.7595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3418 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.898 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 148.225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 642.715 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt2_in[4]
  PIN prt2_in[3] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3916 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.64 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.08 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3816 LAYER M4 ; 
    ANTENNAMAXAREACAR 8.48218 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 11.9754 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA4 ;
  END prt2_in[3]
  PIN prt2_in[2] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 30.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 132.845 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 903.833 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3969.24 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt2_in[2]
  PIN prt2_in[1] 
    ANTENNAPARTIALMETALAREA 0.931 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0964 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 20.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.8368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0451 LAYER M3 ; 
    ANTENNAMAXAREACAR 479.446 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2108.48 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.886918 LAYER VIA3 ;
  END prt2_in[1]
  PIN prt2_in[0] 
    ANTENNAPARTIALMETALAREA 0.5575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.497 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.38679 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 14.6436 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.104822 LAYER VIA2 ;
  END prt2_in[0]
  PIN prt2_out[7] 
    ANTENNAPARTIALMETALAREA 0.471 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0724 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.582 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.2048 LAYER M3 ;
  END prt2_out[7]
  PIN prt2_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.721 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2 ;
  END prt2_out[6]
  PIN prt2_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.759 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4276 LAYER M2 ;
  END prt2_out[5]
  PIN prt2_out[4] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2 ;
  END prt2_out[4]
  PIN prt2_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.521 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3364 LAYER M2 ;
  END prt2_out[3]
  PIN prt2_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.783 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5332 LAYER M2 ;
  END prt2_out[2]
  PIN prt2_out[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.279 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2276 LAYER M2 ;
  END prt2_out[1]
  PIN prt2_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2 ;
  END prt2_out[0]
  PIN prt2_dir[7] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4635 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0394 LAYER M2 ;
  END prt2_dir[7]
  PIN prt2_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2538 LAYER M2 ;
  END prt2_dir[6]
  PIN prt2_dir[5] 
    ANTENNAPARTIALMETALAREA 0.1315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.2608 LAYER M3 ;
  END prt2_dir[5]
  PIN prt2_dir[4] 
    ANTENNAPARTIALMETALAREA 0.3715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6346 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.706 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.1504 LAYER M3 ;
  END prt2_dir[4]
  PIN prt2_dir[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3166 LAYER M2 ;
  END prt2_dir[3]
  PIN prt2_dir[2] 
    ANTENNAPARTIALMETALAREA 0.4135 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8634 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.642 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.0688 LAYER M3 ;
  END prt2_dir[2]
  PIN prt2_dir[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3765 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6566 LAYER M2 ;
  END prt2_dir[1]
  PIN prt2_dir[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2254 LAYER M2 ;
  END prt2_dir[0]
  PIN prt2_ren[7] 
    ANTENNAPARTIALMETALAREA 0.7035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.3008 LAYER M3 ;
  END prt2_ren[7]
  PIN prt2_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5435 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4794 LAYER M2 ;
  END prt2_ren[6]
  PIN prt2_ren[5] 
    ANTENNAPARTIALMETALAREA 0.6945 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0558 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.7808 LAYER M3 ;
  END prt2_ren[5]
  PIN prt2_ren[4] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.9168 LAYER M3 ;
  END prt2_ren[4]
  PIN prt2_ren[3] 
    ANTENNAPARTIALMETALAREA 0.4855 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1802 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.146 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2864 LAYER M3 ;
  END prt2_ren[3]
  PIN prt2_ren[2] 
    ANTENNAPARTIALMETALAREA 0.6675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.937 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.586 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4224 LAYER M3 ;
  END prt2_ren[2]
  PIN prt2_ren[1] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.878 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5072 LAYER M3 ;
  END prt2_ren[1]
  PIN prt2_ren[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3095 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4058 LAYER M2 ;
  END prt2_ren[0]
  PIN prt3_in[7] 
    ANTENNAPARTIALMETALAREA 18.5395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 81.6618 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 537.19 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2364.1 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END prt3_in[7]
  PIN prt3_in[6] 
    ANTENNAPARTIALMETALAREA 15.4885 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 68.2374 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M2 ; 
    ANTENNAMAXAREACAR 573.146 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2523.63 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.369004 LAYER VIA2 ;
  END prt3_in[6]
  PIN prt3_in[5] 
    ANTENNAPARTIALMETALAREA 2.4905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.0022 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 18.228 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.2912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M3 ; 
    ANTENNAMAXAREACAR 632.791 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2787.4 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 1.89702 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.262 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5968 LAYER M4 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 644.949 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 2841.32 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.89702 LAYER VIA4 ;
  END prt3_in[5]
  PIN prt3_in[4] 
    ANTENNAPARTIALMETALAREA 0.2925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.287 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 14.706 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 64.7504 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M5 ; 
    ANTENNAMAXAREACAR 150.916 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 666.035 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.19836 LAYER VIA5 ;
  END prt3_in[4]
  PIN prt3_in[3] 
    ANTENNAPARTIALMETALAREA 0.1755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7722 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 19.19 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.568 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 LAYER M3 ; 
    ANTENNAMAXAREACAR 129.056 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 568.651 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA3 ;
  END prt3_in[3]
  PIN prt3_in[2] 
    ANTENNAPARTIALMETALAREA 2.0335 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9914 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 471.504 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2078.03 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3 ;
  END prt3_in[2]
  PIN prt3_in[1] 
    ANTENNAPARTIALMETALAREA 14.5315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 64.0266 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.7792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 459.769 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2024.77 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3 ;
  END prt3_in[1]
  PIN prt3_in[0] 
    ANTENNAPARTIALMETALAREA 1.8505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1862 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.7488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 409.205 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1783.97 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt3_in[0]
  PIN prt3_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.903 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.6612 LAYER M2 ;
  END prt3_out[7]
  PIN prt3_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.016 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.5584 LAYER M2 ;
  END prt3_out[6]
  PIN prt3_out[5] 
    ANTENNAPARTIALMETALAREA 1.036 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5584 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.726 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6384 LAYER M3 ;
  END prt3_out[5]
  PIN prt3_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.137 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6468 LAYER M2 ;
  END prt3_out[4]
  PIN prt3_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.615 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.394 LAYER M2 ;
  END prt3_out[3]
  PIN prt3_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 9.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 41.448 LAYER M2 ;
  END prt3_out[2]
  PIN prt3_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.25 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.344 LAYER M2 ;
  END prt3_out[1]
  PIN prt3_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.959 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.5076 LAYER M2 ;
  END prt3_out[0]
  PIN prt3_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.8995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.2458 LAYER M2 ;
  END prt3_dir[7]
  PIN prt3_dir[6] 
    ANTENNAPARTIALMETALAREA 5.3565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.5686 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.786 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5024 LAYER M3 ;
  END prt3_dir[6]
  PIN prt3_dir[5] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.206 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M3 ;
  END prt3_dir[5]
  PIN prt3_dir[4] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 15.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 68.5168 LAYER M3 ;
  END prt3_dir[4]
  PIN prt3_dir[3] 
    ANTENNAPARTIALMETALAREA 0.7515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3066 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 16.766 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.8144 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.878 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9072 LAYER M4 ;
  END prt3_dir[3]
  PIN prt3_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.7965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.1486 LAYER M2 ;
  END prt3_dir[2]
  PIN prt3_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.9165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.3646 LAYER M2 ;
  END prt3_dir[1]
  PIN prt3_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.8975 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.881 LAYER M2 ;
  END prt3_dir[0]
  PIN prt3_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.2215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 62.7066 LAYER M2 ;
  END prt3_ren[7]
  PIN prt3_ren[6] 
    ANTENNAPARTIALMETALAREA 4.6185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.3654 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.166 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1744 LAYER M3 ;
  END prt3_ren[6]
  PIN prt3_ren[5] 
    ANTENNAPARTIALMETALAREA 7.3605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.3862 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.042 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.0288 LAYER M3 ;
  END prt3_ren[5]
  PIN prt3_ren[4] 
    ANTENNAPARTIALMETALAREA 0.4005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7622 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.898 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.3952 LAYER M3 ;
  END prt3_ren[4]
  PIN prt3_ren[3] 
    ANTENNAPARTIALMETALAREA 0.2075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.913 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.412 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.3008 LAYER M3 ;
  END prt3_ren[3]
  PIN prt3_ren[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 7.1125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.427 LAYER M2 ;
  END prt3_ren[2]
  PIN prt3_ren[1] 
    ANTENNAPARTIALMETALAREA 11.1805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.1942 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8704 LAYER M3 ;
  END prt3_ren[1]
  PIN prt3_ren[0] 
    ANTENNAPARTIALMETALAREA 0.5805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5542 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.048 LAYER M3 ;
  END prt3_ren[0]
  PIN prt4_in[7] 
    ANTENNAPARTIALMETALAREA 1.3555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9642 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 25.812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 113.661 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 412.374 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1807.8 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.16802 LAYER VIA3 ;
  END prt4_in[7]
  PIN prt4_in[6] 
    ANTENNAPARTIALMETALAREA 1.9355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5162 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 17.758 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.1792 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 5.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.3872 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 67.1771 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 296.923 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA4 ;
  END prt4_in[6]
  PIN prt4_in[5] 
    ANTENNAPARTIALMETALAREA 2.5555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 7.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.4928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.818 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.4432 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 51.23 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 227.415 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.54769 LAYER VIA4 ;
  END prt4_in[5]
  PIN prt4_in[4] 
    ANTENNAPARTIALMETALAREA 6.7775 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.865 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M2 ; 
    ANTENNAMAXAREACAR 184.919 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 814.374 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.813008 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.186 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M3 ;
    ANTENNAGATEAREA 0.0369 LAYER M3 ; 
    ANTENNAMAXAREACAR 189.959 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 837.745 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.622 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7808 LAYER M4 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 195.952 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 864.535 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA4 ;
  END prt4_in[4]
  PIN prt4_in[3] 
    ANTENNAPARTIALMETALAREA 7.2485 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.9814 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M2 ; 
    ANTENNAMAXAREACAR 203.121 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 892.851 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 206.069 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 906.246 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
  END prt4_in[3]
  PIN prt4_in[2] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 290.29 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1277.85 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.62602 LAYER VIA3 ;
  END prt4_in[2]
  PIN prt4_in[1] 
    ANTENNAPARTIALMETALAREA 0.731 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 20.698 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.1152 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 29.0752 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 76.013 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 332.508 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.927362 LAYER VIA4 ;
  END prt4_in[1]
  PIN prt4_in[0] 
    ANTENNAPARTIALMETALAREA 0.2725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 27.886 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 122.742 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 1077.86 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4725.82 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt4_in[0]
  PIN prt4_out[7] 
    ANTENNAPARTIALMETALAREA 10.652 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.7766 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 47.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 52.536 LAYER M3 ;
  END prt4_out[7]
  PIN prt4_out[6] 
    ANTENNAPARTIALMETALAREA 8.572 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4886 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.264 LAYER M3 ;
  END prt4_out[6]
  PIN prt4_out[5] 
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.4902 LAYER M3 ;
  END prt4_out[5]
  PIN prt4_out[4] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5142 LAYER M3 ;
  END prt4_out[4]
  PIN prt4_out[3] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.038 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.6112 LAYER M3 ;
  END prt4_out[3]
  PIN prt4_out[2] 
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.1488 LAYER M3 ;
  END prt4_out[2]
  PIN prt4_out[1] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[1]
  PIN prt4_out[0] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[0]
  PIN prt4_dir[7] 
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.106 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.3104 LAYER M3 ;
  END prt4_dir[7]
  PIN prt4_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2286 LAYER M2 ;
  END prt4_dir[6]
  PIN prt4_dir[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3222 LAYER M2 ;
  END prt4_dir[5]
  PIN prt4_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.4995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5978 LAYER M2 ;
  END prt4_dir[4]
  PIN prt4_dir[3] 
    ANTENNAPARTIALMETALAREA 0.871 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.898 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5952 LAYER M3 ;
  END prt4_dir[3]
  PIN prt4_dir[2] 
    ANTENNAPARTIALMETALAREA 0.491 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1604 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.5408 LAYER M3 ;
  END prt4_dir[2]
  PIN prt4_dir[1] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.722 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.6208 LAYER M6 ;
  END prt4_dir[1]
  PIN prt4_dir[0] 
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6 ;
  END prt4_dir[0]
  PIN prt4_ren[7] 
    ANTENNAPARTIALMETALAREA 0.5075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.233 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.1568 LAYER M3 ;
  END prt4_ren[7]
  PIN prt4_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0534 LAYER M2 ;
  END prt4_ren[6]
  PIN prt4_ren[5] 
    ANTENNAPARTIALMETALAREA 1.2305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4142 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.4368 LAYER M3 ;
  END prt4_ren[5]
  PIN prt4_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.7205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5702 LAYER M2 ;
  END prt4_ren[4]
  PIN prt4_ren[3] 
    ANTENNAPARTIALMETALAREA 3.9985 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6374 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M3 ;
  END prt4_ren[3]
  PIN prt4_ren[2] 
    ANTENNAPARTIALMETALAREA 0.6635 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9194 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.6928 LAYER M3 ;
  END prt4_ren[2]
  PIN prt4_ren[1] 
    ANTENNAPARTIALMETALAREA 0.8035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6 ;
  END prt4_ren[1]
  PIN prt4_ren[0] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.762 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.7968 LAYER M6 ;
  END prt4_ren[0]
  PIN use_dac_glb_bias 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.223 LAYER M2 ;
  END use_dac_glb_bias
  PIN en_bias_buf 
    ANTENNAPARTIALMETALAREA 0.076 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.458 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0592 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.562 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 24.5168 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.078 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 48.7872 LAYER M6 ;
  END en_bias_buf
  PIN en_bias_gen 
    ANTENNAPARTIALMETALAREA 1.839 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1356 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.106 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4032 LAYER M4 ;
  END en_bias_gen
  PIN BIAS_ADJ[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.843 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1972 LAYER M2 ;
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.146 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6864 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.276 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.3024 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M7 ; 
    ANTENNAMAXAREACAR 171.894 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 758.69 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.7316 LAYER VIA7 ;
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.998 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6352 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.818 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 43.2432 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 263.101 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1161.46 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.002 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4528 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.158 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.186 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.6624 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.058 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 48.6992 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 254.301 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1122.74 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.33333 LAYER VIA6 ;
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1] 
    ANTENNAPARTIALMETALAREA 0.122 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5368 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.422 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.718 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.0032 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.996 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 44.0704 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 242.482 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1070.52 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA6 ;
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.678 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4272 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.796 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 43.1904 LAYER M6 ;
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.142 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.922 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7008 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.798 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 47.5552 LAYER M6 ;
  END BIAS_DBP[13]
  PIN BIAS_DBP[12] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.166 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.7744 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 12.9 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 56.848 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 311.957 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1376.05 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6 ;
  END BIAS_DBP[12]
  PIN BIAS_DBP[11] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0816 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.566 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 24.5344 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.698 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 51.5152 LAYER M6 ;
  END BIAS_DBP[11]
  PIN BIAS_DBP[10] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1562 LAYER M2 ;
  END BIAS_DBP[10]
  PIN BIAS_DBP[9] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.002 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.0528 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.576 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 51.0224 LAYER M6 ;
  END BIAS_DBP[9]
  PIN BIAS_DBP[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.341 LAYER M2 ;
  END BIAS_DBP[8]
  PIN BIAS_DBP[7] 
    ANTENNAPARTIALMETALAREA 0.847 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7268 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3568 LAYER M3 ;
  END BIAS_DBP[7]
  PIN BIAS_DBP[6] 
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.164 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.6096 LAYER M3 ;
  END BIAS_DBP[6]
  PIN BIAS_DBP[5] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.456 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 19.6944 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ; 
    ANTENNAMAXAREACAR 141.834 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 630.918 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.18579 LAYER VIA6 ;
  END BIAS_DBP[5]
  PIN BIAS_DBP[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9414 LAYER M2 ;
  END BIAS_DBP[4]
  PIN BIAS_DBP[3] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.062 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3168 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.22 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.656 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.586 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0224 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.92 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 308.184 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1362.93 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_DBP[3]
  PIN BIAS_DBP[2] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.216 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 27.4384 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 240.482 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1065.04 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_DBP[2]
  PIN BIAS_DBP[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
  END BIAS_DBP[1]
  PIN BIAS_DBP[0] 
    ANTENNAPARTIALMETALAREA 0.0885 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.856 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6544 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.726 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.0384 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.578 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 24.5872 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 211.828 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 935.061 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6 ;
  END BIAS_DBP[0]
  PIN BIAS_DBN[13] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.958 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.498 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6352 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.338 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9312 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.364 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 32.4896 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 119.773 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 529.356 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_DBN[13]
  PIN BIAS_DBN[12] 
    ANTENNAPARTIALMETALAREA 1.4055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1842 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.086 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4224 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.968 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.738 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 20.8912 LAYER M6 ;
  END BIAS_DBN[12]
  PIN BIAS_DBN[11] 
    ANTENNAPARTIALMETALAREA 2.597 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4268 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.968 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.002 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6528 LAYER M4 ;
  END BIAS_DBN[11]
  PIN BIAS_DBN[10] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.968 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.538 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.4112 LAYER M4 ;
  END BIAS_DBN[10]
  PIN BIAS_DBN[9] 
    ANTENNAPARTIALMETALAREA 0.05 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER M3 ;
  END BIAS_DBN[9]
  PIN BIAS_DBN[8] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.678 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0272 LAYER M4 ;
  END BIAS_DBN[8]
  PIN BIAS_DBN[7] 
    ANTENNAPARTIALMETALAREA 0.513 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3012 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.138 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M3 ;
  END BIAS_DBN[7]
  PIN BIAS_DBN[6] 
    ANTENNAPARTIALMETALAREA 0.4515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0306 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.158 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M3 ;
  END BIAS_DBN[6]
  PIN BIAS_DBN[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.962 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.978 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.246 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.518 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 28.7232 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 356.214 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1572.49 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_DBN[5]
  PIN BIAS_DBN[4] 
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.498 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.0352 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.506 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2704 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.278 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 32.0672 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER M6 ; 
    ANTENNAMAXAREACAR 163.191 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 721.322 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.4245 LAYER VIA6 ;
  END BIAS_DBN[4]
  PIN BIAS_DBN[3] 
    ANTENNAPARTIALMETALAREA 0.833 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6652 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.766 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4144 LAYER M3 ;
  END BIAS_DBN[3]
  PIN BIAS_DBN[2] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.282 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.2848 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.404 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 41.4656 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 210.85 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 929.492 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA6 ;
  END BIAS_DBN[2]
  PIN BIAS_DBN[1] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.362 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.2368 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.874 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.7776 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 444.305 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1960.55 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_DBN[1]
  PIN BIAS_DBN[0] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.698 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1152 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.962 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6768 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.098 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.0752 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 260.281 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1148.84 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6 ;
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13] 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.71 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.212 LAYER M2 ;
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4322 LAYER M2 ;
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2882 LAYER M2 ;
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0684 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.044 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 26.6816 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 4.642 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.4688 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.622 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 33.5808 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 393.568 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1734.15 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA6 ;
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.506 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 13.234 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 58.3616 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 2.938 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0592 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 168.973 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 747.939 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA7 ;
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.958 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6592 LAYER M4 ;
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.748 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3792 LAYER M3 ;
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3] 
    ANTENNAPARTIALMETALAREA 0.142 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6248 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.548 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER M3 ;
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2] 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.818 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 30.0432 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 254.402 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1119.75 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA4 ;
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1] 
    ANTENNAPARTIALMETALAREA 0.051 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2244 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7808 LAYER M3 ;
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0] 
    ANTENNAPARTIALMETALAREA 0.2445 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1198 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.3168 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2512 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.832 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.5928 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.564 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 20.1696 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 25.2836 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 114.411 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.77994 LAYER VIA7 ;
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.318 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.6432 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.922 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7008 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.062 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7168 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.522 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 19.9408 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 134.417 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 595.688 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12] 
    ANTENNAPARTIALMETALAREA 0.502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1264 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.478 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.9472 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.086 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4224 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.338 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.5312 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 123.299 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 546.133 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11] 
    ANTENNAPARTIALMETALAREA 0.358 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6192 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.878 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7072 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.968 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.538 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6112 LAYER M6 ;
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 3.018 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3232 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.198 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 27.3152 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 96.1201 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 425.911 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA6 ;
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.422 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.226 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.118 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.1632 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 185.368 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 818.703 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA6 ;
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8] 
    ANTENNAPARTIALMETALAREA 0.1415 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.618 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 29.1632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 2.618 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5632 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 105.601 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 467.73 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7] 
    ANTENNAPARTIALMETALAREA 0.102 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4488 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.858 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 34.6192 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.302 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M5 ; 
    ANTENNAMAXAREACAR 21.3408 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 90.5033 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA5 ;
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.418 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8832 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 7.176 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 31.6624 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 0.126 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M7 ; 
    ANTENNAMAXAREACAR 22.9342 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 104.73 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.83333 LAYER VIA7 ;
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.326 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4784 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.142 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.3568 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 464.871 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2053.54 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4] 
    ANTENNAPARTIALMETALAREA 0.0215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0946 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M3 ;
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.978 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 30.7472 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 LAYER M6 ; 
    ANTENNAMAXAREACAR 187.406 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 815.547 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.64609 LAYER VIA6 ;
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2] 
    ANTENNAPARTIALMETALAREA 0.0545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.982 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3648 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.158 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7392 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.386 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5424 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.318 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 32.2432 LAYER M6 ;
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1] 
    ANTENNAPARTIALMETALAREA 0.023 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1012 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5648 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4112 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.742 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7088 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.916 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 30.5184 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 0.126 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M7 ; 
    ANTENNAMAXAREACAR 177.686 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 788.505 LAYER M7 ;
    ANTENNAMAXCUTCAR 3.55987 LAYER VIA7 ;
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0] 
    ANTENNAPARTIALMETALAREA 0.0195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.478 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1472 LAYER M4 ;
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.131 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.4835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1714 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.8592 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 53.0667 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4] 
    ANTENNAPARTIALMETALAREA 1.043 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.96 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 15.1 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 66.528 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.282 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 5.392 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 23.8128 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0411 LAYER M7 ; 
    ANTENNAMAXAREACAR 782.012 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 3436.03 LAYER M7 ;
    ANTENNAMAXCUTCAR 2.91971 LAYER VIA7 ;
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.6165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.493 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2132 LAYER M2 ;
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.3505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5422 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.758 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.3916 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 152.317 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.323625 LAYER VIA3 ;
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.241 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4604 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M2 ; 
    ANTENNAMAXAREACAR 20.8803 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 91.4434 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.161812 LAYER VIA2 ;
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.2505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1022 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.488 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.0352 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 44.7167 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 198.403 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4] 
    ANTENNAPARTIALMETALAREA 0.224 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9856 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.802 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5728 LAYER M3 ;
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.087 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3828 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.4995 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2418 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.526 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 43.7167 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 194.737 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA4 ;
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.782 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.6833 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.323 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.1375 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.605 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.338 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9312 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 62.2091 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 274.036 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA4 ;
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7432 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.978 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.4009 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 77.3204 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.323625 LAYER VIA3 ;
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[15] 
    ANTENNAPARTIALMETALAREA 0.1335 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5874 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 4.396 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.4304 LAYER M5 ;
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14] 
    ANTENNAPARTIALMETALAREA 0.511 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2484 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.486 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1824 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 7.118 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 31.3632 LAYER M5 ;
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13] 
    ANTENNAPARTIALMETALAREA 0.4695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0658 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.5808 LAYER M3 ;
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12] 
    ANTENNAPARTIALMETALAREA 0.331 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.1792 LAYER M3 ;
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11] 
    ANTENNAPARTIALMETALAREA 0.071 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3124 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.438 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7712 LAYER M5 ;
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10] 
    ANTENNAPARTIALMETALAREA 0.249 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0956 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.6848 LAYER M3 ;
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.342 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M2 ;
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8] 
    ANTENNAPARTIALMETALAREA 0.075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.33 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.624 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0336 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.206 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M6 ;
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5295 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3298 LAYER M2 ;
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6] 
    ANTENNAPARTIALMETALAREA 1.287 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.788 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3552 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.586 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 24.158 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 106.339 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.102 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 2.602 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4928 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0481 LAYER M7 ; 
    ANTENNAMAXAREACAR 279.371 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 1235.97 LAYER M7 ;
    ANTENNAMAXCUTCAR 2.2869 LAYER VIA7 ;
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4145 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8678 LAYER M2 ;
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.466 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0944 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6992 LAYER M4 ;
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3] 
    ANTENNAPARTIALMETALAREA 0.431 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8964 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.3785 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1094 LAYER M3 ;
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.29 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32 LAYER M2 ;
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1] 
    ANTENNAPARTIALMETALAREA 0.0915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4026 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9488 LAYER M3 ;
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0] 
    ANTENNAPARTIALMETALAREA 0.154 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4032 LAYER M4 ;
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0752 LAYER M4 ;
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.378 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1072 LAYER M4 ;
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3088 LAYER M3 ;
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6992 LAYER M4 ;
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.358 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3752 LAYER M2 ;
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.3705 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0742 LAYER M2 ;
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.106 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M2 ;
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.906 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0304 LAYER M3 ;
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.217 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9988 LAYER M2 ;
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4] 
    ANTENNAPARTIALMETALAREA 0.0305 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1342 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M3 ;
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3] 
    ANTENNAPARTIALMETALAREA 0.068 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.726 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2384 LAYER M3 ;
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2] 
    ANTENNAPARTIALMETALAREA 0.0195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.818 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6432 LAYER M3 ;
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1] 
    ANTENNAPARTIALMETALAREA 0.074 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3256 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.782 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4848 LAYER M3 ;
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4158 LAYER M2 ;
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.5375 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.409 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.87374 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 42.2165 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.6544 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.4863 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.978 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3472 LAYER M4 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 27.767 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 122.216 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.865801 LAYER VIA4 ;
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.498 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.9912 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 29.816 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 131.278 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.166 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 27.1744 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M6 ; 
    ANTENNAMAXAREACAR 390.539 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1721.21 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA6 ;
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2902 LAYER M2 ;
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 1.379 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0676 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M2 ; 
    ANTENNAMAXAREACAR 20.8189 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 90.3867 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.446 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0064 LAYER M3 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.2547 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.339 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.4329 LAYER VIA3 ;
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.7975 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.509 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.886 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9424 LAYER M3 ;
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9512 LAYER M2 ;
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.1115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4906 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.658 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9392 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 122.506 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 538.984 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA4 ;
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.551 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4244 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.432 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.582 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6048 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.558 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 49.4664 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 214.252 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA5 ;
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.1225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.1424 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7696 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.218 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2032 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 64.3912 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 285.502 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA5 ;
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.047 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.142 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0688 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.942 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9888 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 79.0376 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 347.744 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA5 ;
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.1775 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.781 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.366 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6544 LAYER M3 ;
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.391 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7204 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M3 ;
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4885 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1494 LAYER M2 ;
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4] 
    ANTENNAPARTIALMETALAREA 1.107 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8708 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.896 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.8304 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.9806 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 217.107 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.371 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.138 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.1 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.928 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.286 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1024 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 55.6214 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 247.152 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA5 ;
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.129 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5676 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.958 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 79.1489 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 349.961 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.809061 LAYER VIA4 ;
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.1665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.685 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.014 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.438 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9712 LAYER M3 ;
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.7015 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0866 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.858 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8192 LAYER M3 ;
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.696 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.19 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ; 
    ANTENNAMAXAREACAR 95.7067 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 421.249 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.666667 LAYER VIA3 ;
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.553 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4772 LAYER M2 ;
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.694 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.898 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9952 LAYER M3 ;
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.6195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7258 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.418 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2832 LAYER M3 ;
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5 LAYER M2 ;
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.993 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.0572 LAYER M2 ;
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.698 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1152 LAYER M4 ;
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11] 
    ANTENNAPARTIALMETALAREA 0.05 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.948 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M3 ;
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.122 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5808 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6672 LAYER M4 ;
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.818 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6432 LAYER M4 ;
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.142 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M3 ;
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8048 LAYER M3 ;
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6] 
    ANTENNAPARTIALMETALAREA 0.0185 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.344 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6016 LAYER M2 ;
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.3295 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4938 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.298 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7552 LAYER M4 ;
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7808 LAYER M3 ;
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.308 LAYER M2 ;
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.165 LAYER M2 ;
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done 
    ANTENNAPARTIALMETALAREA 0.186 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.142 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.8688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 341.62 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1504.42 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.755668 LAYER VIA3 ;
  END dsadc_conv_done
  PIN dsadc_en 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.237 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0868 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.682 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0448 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.804 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 25.6256 LAYER M5 ;
  END dsadc_en
  PIN dsadc_clk 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.224 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3224 LAYER M3 ;
  END dsadc_clk
  PIN dsadc_switch[2] 
    ANTENNAPARTIALMETALAREA 0.111 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4884 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.1205 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5742 LAYER M3 ;
  END dsadc_switch[2]
  PIN dsadc_switch[1] 
    ANTENNAPARTIALMETALAREA 0.584 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5696 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.618 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1632 LAYER M3 ;
  END dsadc_switch[1]
  PIN dsadc_switch[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.291 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2804 LAYER M2 ;
  END dsadc_switch[0]
  PIN dac_en_pot 
    ANTENNAPARTIALMETALAREA 0.1665 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.198 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.9152 LAYER M5 ;
  END dac_en_pot
  PIN adc_ext_in 
    ANTENNAPARTIALMETALAREA 0.571 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5124 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.198 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.5152 LAYER M3 ;
  END adc_ext_in
  PIN atp_en 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.562 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5168 LAYER M4 ;
  END atp_en
  PIN atp_sel 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.364 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6456 LAYER M2 ;
  END atp_sel
  PIN adc_sel 
    ANTENNAPARTIALMETALAREA 0.3095 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.922 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.3008 LAYER M3 ;
  END adc_sel
  PIN saradc_clk 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 65.902 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 72.6682 LAYER M3 ;
  END saradc_clk
  PIN saradc_rdy 
    ANTENNAPARTIALMETALAREA 0.481 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2484 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 25.5908 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 110.807 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END saradc_rdy
  PIN saradc_rst 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.291 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2804 LAYER M2 ;
  END saradc_rst
  PIN saradc_data[9] 
    ANTENNAPARTIALMETALAREA 0.8825 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.883 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.4128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 272.166 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1190.89 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END saradc_data[9]
  PIN saradc_data[8] 
    ANTENNAPARTIALMETALAREA 0.4055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8282 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 6.378 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.1072 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M4 ; 
    ANTENNAMAXAREACAR 47.5642 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 211.683 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.25945 LAYER VIA4 ;
  END saradc_data[8]
  PIN saradc_data[7] 
    ANTENNAPARTIALMETALAREA 0.4315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.1648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 279.37 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1226.55 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END saradc_data[7]
  PIN saradc_data[6] 
    ANTENNAPARTIALMETALAREA 0.271 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.1335 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.0314 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 290.249 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1267.37 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END saradc_data[6]
  PIN saradc_data[5] 
    ANTENNAPARTIALMETALAREA 0.6755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9722 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.098 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8752 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.266 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 12.638 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 55.6512 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 1.358 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0192 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M6 ; 
    ANTENNAMAXAREACAR 125.013 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 547.259 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.51889 LAYER VIA6 ;
  END saradc_data[5]
  PIN saradc_data[4] 
    ANTENNAPARTIALMETALAREA 0.5465 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4046 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 9.158 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.3392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 246.725 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1083.64 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END saradc_data[4]
  PIN saradc_data[3] 
    ANTENNAPARTIALMETALAREA 0.1825 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.803 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 9.818 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 43.2432 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5 ; 
    ANTENNAMAXAREACAR 342.393 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1508.99 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.01511 LAYER VIA5 ;
  END saradc_data[3]
  PIN saradc_data[2] 
    ANTENNAPARTIALMETALAREA 0.6425 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.827 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.5792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M3 ; 
    ANTENNAMAXAREACAR 304.861 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1338.35 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.00756 LAYER VIA3 ;
  END saradc_data[2]
  PIN saradc_data[1] 
    ANTENNAPARTIALMETALAREA 0.171 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7524 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.3135 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8234 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.606 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7104 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 9.938 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 43.7712 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5 ; 
    ANTENNAMAXAREACAR 390.453 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1721.18 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.01511 LAYER VIA5 ;
  END saradc_data[1]
  PIN saradc_data[0] 
    ANTENNAPARTIALMETALAREA 0.0395 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1738 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.566 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.678 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 60.2272 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0397 LAYER M5 ; 
    ANTENNAMAXAREACAR 419.27 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1846.5 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.76322 LAYER VIA5 ;
  END saradc_data[0]
END MCU

END LIBRARY
