

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO MCU 
  PIN resetn_in 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 25.802 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 113.573 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M6 ; 
    ANTENNAMAXAREACAR 973.496 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4290.04 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.32103 LAYER VIA6 ;
  END resetn_in
  PIN resetn_out 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.474 LAYER M2 ;
  END resetn_out
  PIN resetn_dir 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6365 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8446 LAYER M2 ;
  END resetn_dir
  PIN resetn_ren 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5895 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6378 LAYER M2 ;
  END resetn_ren
  PIN prt1_in[7] 
    ANTENNAPARTIALMETALAREA 4.0155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6682 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 11.398 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.1952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 357.85 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1556.14 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt1_in[7]
  PIN prt1_in[6] 
    ANTENNAPARTIALMETALAREA 22.8945 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 100.78 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.5808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 128.484 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 556.133 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA3 ;
  END prt1_in[6]
  PIN prt1_in[5] 
    ANTENNAPARTIALMETALAREA 0.0725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.319 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 14.456 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.6944 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2577 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.2742 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 264.591 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.467722 LAYER VIA3 ;
  END prt1_in[5]
  PIN prt1_in[4] 
    ANTENNAPARTIALMETALAREA 5.5325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.343 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 14.692 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.7328 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2577 LAYER M3 ; 
    ANTENNAMAXAREACAR 63.5292 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 279.233 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.747384 LAYER VIA3 ;
  END prt1_in[4]
  PIN prt1_in[3] 
    ANTENNAPARTIALMETALAREA 0.496 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5456 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4982 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.65068 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.9518 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.314465 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4422 LAYER M4 ;
    ANTENNAGATEAREA 0.1908 LAYER M4 ; 
    ANTENNAMAXAREACAR 10.919 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 19.2694 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 0.419287 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.28 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER M5 ;
    ANTENNAGATEAREA 0.2544 LAYER M5 ; 
    ANTENNAMAXAREACAR 21.8821 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 36.2516 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.10063 LAYER VIA5 ;
  END prt1_in[3]
  PIN prt1_in[2] 
    ANTENNAPARTIALMETALAREA 6.3935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.1754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 6.246 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.5264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 87.7248 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 385.805 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[2]
  PIN prt1_in[1] 
    ANTENNAPARTIALMETALAREA 14.6155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 64.3082 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 8.806 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.7904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M3 ; 
    ANTENNAMAXAREACAR 114.772 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 500.057 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.453001 LAYER VIA3 ;
  END prt1_in[1]
  PIN prt1_in[0] 
    ANTENNAPARTIALMETALAREA 1.3755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0522 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.718 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.0032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0447 LAYER M3 ; 
    ANTENNAMAXAREACAR 424.193 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1868.05 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.671141 LAYER VIA3 ;
  END prt1_in[0]
  PIN prt1_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 7.418 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.6832 LAYER M2 ;
  END prt1_out[7]
  PIN prt1_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.179 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.0756 LAYER M2 ;
  END prt1_out[6]
  PIN prt1_out[5] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[5]
  PIN prt1_out[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[4]
  PIN prt1_out[3] 
    ANTENNAPARTIALMETALAREA 0.976 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2944 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.726 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.8384 LAYER M3 ;
  END prt1_out[3]
  PIN prt1_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[2]
  PIN prt1_out[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2948 LAYER M2 ;
  END prt1_out[1]
  PIN prt1_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.255 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.61 LAYER M2 ;
  END prt1_out[0]
  PIN prt1_dir[7] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[7]
  PIN prt1_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.7595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.2298 LAYER M2 ;
  END prt1_dir[6]
  PIN prt1_dir[5] 
    ANTENNAPARTIALMETALAREA 4.9005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5622 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.2992 LAYER M3 ;
  END prt1_dir[5]
  PIN prt1_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1215 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5786 LAYER M2 ;
  END prt1_dir[4]
  PIN prt1_dir[3] 
    ANTENNAPARTIALMETALAREA 0.5565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.466 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.6944 LAYER M3 ;
  END prt1_dir[3]
  PIN prt1_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5566 LAYER M2 ;
  END prt1_dir[2]
  PIN prt1_dir[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt1_dir[1]
  PIN prt1_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 12.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 53.0926 LAYER M2 ;
  END prt1_dir[0]
  PIN prt1_ren[7] 
    ANTENNAPARTIALMETALAREA 0.1005 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4422 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.466 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4944 LAYER M3 ;
  END prt1_ren[7]
  PIN prt1_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.4235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.1514 LAYER M2 ;
  END prt1_ren[6]
  PIN prt1_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.9835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 66.0154 LAYER M2 ;
  END prt1_ren[5]
  PIN prt1_ren[4] 
    ANTENNAPARTIALMETALAREA 4.2225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.623 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.6208 LAYER M3 ;
  END prt1_ren[4]
  PIN prt1_ren[3] 
    ANTENNAPARTIALMETALAREA 0.2475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.089 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.586 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8224 LAYER M3 ;
  END prt1_ren[3]
  PIN prt1_ren[2] 
    ANTENNAPARTIALMETALAREA 1.5455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.732 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5088 LAYER M3 ;
  END prt1_ren[2]
  PIN prt1_ren[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
  END prt1_ren[1]
  PIN prt1_ren[0] 
    ANTENNAPARTIALMETALAREA 0.3675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
  END prt1_ren[0]
  PIN prt2_in[7] 
    ANTENNAPARTIALMETALAREA 0.7535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3594 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0595 LAYER M2 ; 
    ANTENNAMAXAREACAR 15.8361 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 68.6218 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.336134 LAYER VIA2 ;
  END prt2_in[7]
  PIN prt2_in[6] 
    ANTENNAPARTIALMETALAREA 0.4975 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.233 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M2 ; 
    ANTENNAMAXAREACAR 22.9539 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 97.9135 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.576369 LAYER VIA2 ;
  END prt2_in[6]
  PIN prt2_in[5] 
    ANTENNAPARTIALMETALAREA 0.7745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4518 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0883 LAYER M2 ; 
    ANTENNAMAXAREACAR 9.65572 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 41.8029 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.226501 LAYER VIA2 ;
  END prt2_in[5]
  PIN prt2_in[4] 
    ANTENNAPARTIALMETALAREA 0.7955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5002 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 5.642 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.8688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 170.703 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 741.205 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt2_in[4]
  PIN prt2_in[3] 
    ANTENNAPARTIALMETALAREA 0.174 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1914 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.244 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4444 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER M4 ; 
    ANTENNAMAXAREACAR 6.24203 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 8.86751 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.125786 LAYER VIA4 ;
  END prt2_in[3]
  PIN prt2_in[2] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 23.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 103.013 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M3 ; 
    ANTENNAMAXAREACAR 722.334 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3162.55 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15274 LAYER VIA3 ;
  END prt2_in[2]
  PIN prt2_in[1] 
    ANTENNAPARTIALMETALAREA 0.3555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5642 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 15.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.3904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0451 LAYER M3 ; 
    ANTENNAMAXAREACAR 372.262 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1627.45 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.886918 LAYER VIA3 ;
  END prt2_in[1]
  PIN prt2_in[0] 
    ANTENNAPARTIALMETALAREA 0.3535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5994 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.73585 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 15.9135 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.157233 LAYER VIA2 ;
  END prt2_in[0]
  PIN prt2_out[7] 
    ANTENNAPARTIALMETALAREA 0.471 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0724 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.6992 LAYER M3 ;
  END prt2_out[7]
  PIN prt2_out[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.721 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2 ;
  END prt2_out[6]
  PIN prt2_out[5] 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2288 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.378 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7072 LAYER M3 ;
  END prt2_out[5]
  PIN prt2_out[4] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.292 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M2 ;
  END prt2_out[4]
  PIN prt2_out[3] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2 ;
  END prt2_out[3]
  PIN prt2_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.735 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.322 LAYER M2 ;
  END prt2_out[2]
  PIN prt2_out[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.279 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2276 LAYER M2 ;
  END prt2_out[1]
  PIN prt2_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.312 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M2 ;
  END prt2_out[0]
  PIN prt2_dir[7] 
    ANTENNAPARTIALMETALAREA 0.6565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8886 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.1648 LAYER M3 ;
  END prt2_dir[7]
  PIN prt2_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2538 LAYER M2 ;
  END prt2_dir[6]
  PIN prt2_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4254 LAYER M2 ;
  END prt2_dir[5]
  PIN prt2_dir[4] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1946 LAYER M2 ;
  END prt2_dir[4]
  PIN prt2_dir[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3486 LAYER M2 ;
  END prt2_dir[3]
  PIN prt2_dir[2] 
    ANTENNAPARTIALMETALAREA 0.6985 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0734 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.5408 LAYER M3 ;
  END prt2_dir[2]
  PIN prt2_dir[1] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.6835 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0074 LAYER M2 ;
  END prt2_dir[1]
  PIN prt2_dir[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2545 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1198 LAYER M2 ;
  END prt2_dir[0]
  PIN prt2_ren[7] 
    ANTENNAPARTIALMETALAREA 0.7035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.4288 LAYER M3 ;
  END prt2_ren[7]
  PIN prt2_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.7035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1834 LAYER M2 ;
  END prt2_ren[6]
  PIN prt2_ren[5] 
    ANTENNAPARTIALMETALAREA 0.6505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8622 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.642 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2688 LAYER M3 ;
  END prt2_ren[5]
  PIN prt2_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.519 LAYER M2 ;
  END prt2_ren[4]
  PIN prt2_ren[3] 
    ANTENNAPARTIALMETALAREA 0.6675 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.937 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.486 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.1824 LAYER M3 ;
  END prt2_ren[3]
  PIN prt2_ren[2] 
    ANTENNAPARTIALMETALAREA 0.9315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.038 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.4112 LAYER M3 ;
  END prt2_ren[2]
  PIN prt2_ren[1] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2078 LAYER M2 ;
  END prt2_ren[1]
  PIN prt2_ren[0] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4765 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1406 LAYER M2 ;
  END prt2_ren[0]
  PIN prt3_in[7] 
    ANTENNAPARTIALMETALAREA 18.7995 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 82.8058 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M2 ; 
    ANTENNAMAXAREACAR 772.782 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3400.25 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.816327 LAYER VIA2 ;
  END prt3_in[7]
  PIN prt3_in[6] 
    ANTENNAPARTIALMETALAREA 16.2905 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 71.7222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 14.898 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.5952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 569.225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2500.84 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[6]
  PIN prt3_in[5] 
    ANTENNAPARTIALMETALAREA 7.2565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.9286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 14.798 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.1552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 LAYER M3 ; 
    ANTENNAMAXAREACAR 405.474 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1786.01 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.242 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9088 LAYER M4 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 427.073 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1881.47 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.35501 LAYER VIA4 ;
  END prt3_in[5]
  PIN prt3_in[4] 
    ANTENNAPARTIALMETALAREA 0.6325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.783 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.7808 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.178 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8272 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.154 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.7216 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M5 ; 
    ANTENNAMAXAREACAR 76.202 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 337.434 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.16802 LAYER VIA5 ;
  END prt3_in[4]
  PIN prt3_in[3] 
    ANTENNAPARTIALMETALAREA 5.4755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.0922 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 17.934 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.9536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 LAYER M3 ; 
    ANTENNAMAXAREACAR 138.186 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 607.638 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.08401 LAYER VIA3 ;
  END prt3_in[3]
  PIN prt3_in[2] 
    ANTENNAPARTIALMETALAREA 6.1015 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.8906 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 13.538 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.6112 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 542.524 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2361.33 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[2]
  PIN prt3_in[1] 
    ANTENNAPARTIALMETALAREA 14.8155 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.2762 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.9248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 177.269 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 762.155 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt3_in[1]
  PIN prt3_in[0] 
    ANTENNAPARTIALMETALAREA 23.4935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 103.415 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 4.938 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 353.496 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1557.17 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.10701 LAYER VIA3 ;
  END prt3_in[0]
  PIN prt3_out[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.781 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.1684 LAYER M2 ;
  END prt3_out[7]
  PIN prt3_out[6] 
    ANTENNAPARTIALMETALAREA 6.334 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9136 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
  END prt3_out[6]
  PIN prt3_out[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.137 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6468 LAYER M2 ;
  END prt3_out[5]
  PIN prt3_out[4] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.157 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7348 LAYER M2 ;
  END prt3_out[4]
  PIN prt3_out[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3124 LAYER M2 ;
  END prt3_out[3]
  PIN prt3_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 11.337 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.0148 LAYER M2 ;
  END prt3_out[2]
  PIN prt3_out[1] 
    ANTENNAPARTIALMETALAREA 6.816 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.9904 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.484 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.062 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7168 LAYER M4 ;
  END prt3_out[1]
  PIN prt3_out[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.039 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.8596 LAYER M2 ;
  END prt3_out[0]
  PIN prt3_dir[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.9035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.2634 LAYER M2 ;
  END prt3_dir[7]
  PIN prt3_dir[6] 
    ANTENNAPARTIALMETALAREA 5.0385 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.786 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5024 LAYER M3 ;
  END prt3_dir[6]
  PIN prt3_dir[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt3_dir[5]
  PIN prt3_dir[4] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0515 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2266 LAYER M2 ;
  END prt3_dir[4]
  PIN prt3_dir[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER M2 ;
  END prt3_dir[3]
  PIN prt3_dir[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.476 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.3824 LAYER M2 ;
  END prt3_dir[2]
  PIN prt3_dir[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.9745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 61.5758 LAYER M2 ;
  END prt3_dir[1]
  PIN prt3_dir[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.9955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3562 LAYER M2 ;
  END prt3_dir[0]
  PIN prt3_ren[7] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 13.5635 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.7674 LAYER M2 ;
  END prt3_ren[7]
  PIN prt3_ren[6] 
    ANTENNAPARTIALMETALAREA 4.8585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.4214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.026 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3584 LAYER M3 ;
  END prt3_ren[6]
  PIN prt3_ren[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 6.9815 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.8506 LAYER M2 ;
  END prt3_ren[5]
  PIN prt3_ren[4] 
    ANTENNAPARTIALMETALAREA 0.2605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1462 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.758 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.1792 LAYER M3 ;
  END prt3_ren[4]
  PIN prt3_ren[3] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.268 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.0672 LAYER M3 ;
  END prt3_ren[3]
  PIN prt3_ren[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 8.1125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.827 LAYER M2 ;
  END prt3_ren[2]
  PIN prt3_ren[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.3925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 63.459 LAYER M2 ;
  END prt3_ren[1]
  PIN prt3_ren[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 2.4875 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.033 LAYER M2 ;
  END prt3_ren[0]
  PIN prt4_in[7] 
    ANTENNAPARTIALMETALAREA 1.7555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 25.062 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 110.317 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.1872 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 79.9916 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 348.865 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.81869 LAYER VIA4 ;
  END prt4_in[7]
  PIN prt4_in[6] 
    ANTENNAPARTIALMETALAREA 2.9755 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0922 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 17.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M3 ; 
    ANTENNAMAXAREACAR 176.889 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 776.491 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.734684 LAYER VIA3 ;
  END prt4_in[6]
  PIN prt4_in[5] 
    ANTENNAPARTIALMETALAREA 1.6585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2974 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 7.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.438 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7712 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 50.9484 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 224.404 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.927362 LAYER VIA4 ;
  END prt4_in[5]
  PIN prt4_in[4] 
    ANTENNAPARTIALMETALAREA 4.2015 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.5306 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.3509 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 189.742 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.542005 LAYER VIA2 ;
  END prt4_in[4]
  PIN prt4_in[3] 
    ANTENNAPARTIALMETALAREA 0.0525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.438 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.1712 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 6.218 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.4032 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 82.0963 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 362.803 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.00569 LAYER VIA4 ;
  END prt4_in[3]
  PIN prt4_in[2] 
    ANTENNAPARTIALMETALAREA 0.6725 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.959 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 12.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.6448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 5.258 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.1792 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 75.9197 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 335.046 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.81869 LAYER VIA4 ;
  END prt4_in[2]
  PIN prt4_in[1] 
    ANTENNAPARTIALMETALAREA 0.731 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2164 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 20.718 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.2032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 5.858 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.8192 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1038 LAYER M4 ; 
    ANTENNAMAXAREACAR 80.3159 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 353.92 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.734684 LAYER VIA4 ;
  END prt4_in[1]
  PIN prt4_in[0] 
    ANTENNAPARTIALMETALAREA 0.2925 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.287 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 28.622 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 125.981 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M3 ; 
    ANTENNAMAXAREACAR 1087.84 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4765.23 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.47601 LAYER VIA3 ;
  END prt4_in[0]
  PIN prt4_out[7] 
    ANTENNAPARTIALMETALAREA 5.292 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8806 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 81.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.848 LAYER M3 ;
  END prt4_out[7]
  PIN prt4_out[6] 
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 24.562 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.1942 LAYER M3 ;
  END prt4_out[6]
  PIN prt4_out[5] 
    ANTENNAPARTIALMETALAREA 0.172 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1892 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.9142 LAYER M3 ;
  END prt4_out[5]
  PIN prt4_out[4] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.602 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9382 LAYER M3 ;
  END prt4_out[4]
  PIN prt4_out[3] 
    ANTENNAPARTIALMETALAREA 0.831 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6564 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.798 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.5552 LAYER M3 ;
  END prt4_out[3]
  PIN prt4_out[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.719 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2516 LAYER M2 ;
  END prt4_out[2]
  PIN prt4_out[1] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.922 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 74.5008 LAYER M6 ;
  END prt4_out[1]
  PIN prt4_out[0] 
    ANTENNAPARTIALMETALAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5328 LAYER M6 ;
  END prt4_out[0]
  PIN prt4_dir[7] 
    ANTENNAPARTIALMETALAREA 0.631 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7764 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.098 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.2752 LAYER M3 ;
  END prt4_dir[7]
  PIN prt4_dir[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3165 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4366 LAYER M2 ;
  END prt4_dir[6]
  PIN prt4_dir[5] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2765 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2166 LAYER M2 ;
  END prt4_dir[5]
  PIN prt4_dir[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8554 LAYER M2 ;
  END prt4_dir[4]
  PIN prt4_dir[3] 
    ANTENNAPARTIALMETALAREA 0.871 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8324 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.968 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.902 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.6128 LAYER M3 ;
  END prt4_dir[3]
  PIN prt4_dir[2] 
    ANTENNAPARTIALMETALAREA 0.911 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0084 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.338 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.7312 LAYER M3 ;
  END prt4_dir[2]
  PIN prt4_dir[1] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0768 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.722 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.6208 LAYER M6 ;
  END prt4_dir[1]
  PIN prt4_dir[0] 
    ANTENNAPARTIALMETALAREA 0.7795 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4298 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6 ;
  END prt4_dir[0]
  PIN prt4_ren[7] 
    ANTENNAPARTIALMETALAREA 0.5075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.233 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.1568 LAYER M3 ;
  END prt4_ren[7]
  PIN prt4_ren[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.9475 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.257 LAYER M2 ;
  END prt4_ren[6]
  PIN prt4_ren[5] 
    ANTENNAPARTIALMETALAREA 1.0505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.646 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.6864 LAYER M3 ;
  END prt4_ren[5]
  PIN prt4_ren[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.5275 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.721 LAYER M2 ;
  END prt4_ren[4]
  PIN prt4_ren[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1785 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2294 LAYER M2 ;
  END prt4_ren[3]
  PIN prt4_ren[2] 
    ANTENNAPARTIALMETALAREA 0.5035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2154 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.3088 LAYER M3 ;
  END prt4_ren[2]
  PIN prt4_ren[1] 
    ANTENNAPARTIALMETALAREA 0.8035 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 15.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 70.1888 LAYER M6 ;
  END prt4_ren[1]
  PIN prt4_ren[0] 
    ANTENNAPARTIALMETALAREA 0.0405 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1782 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 16.762 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.7968 LAYER M6 ;
  END prt4_ren[0]
  PIN use_dac_glb_bias 
    ANTENNAPARTIALMETALAREA 0.0575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.253 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2512 LAYER M4 ;
  END use_dac_glb_bias
  PIN en_bias_buf 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3124 LAYER M2 ;
  END en_bias_buf
  PIN en_bias_gen 
    ANTENNAPARTIALMETALAREA 0.619 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7676 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.678 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4272 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 4.306 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.9904 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.628 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 46.8512 LAYER M6 ;
  END en_bias_gen
  PIN BIAS_ADJ[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.594 LAYER M2 ;
  END BIAS_ADJ[5]
  PIN BIAS_ADJ[4] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
  END BIAS_ADJ[4]
  PIN BIAS_ADJ[3] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.702 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1328 LAYER M3 ;
  END BIAS_ADJ[3]
  PIN BIAS_ADJ[2] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.546 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8464 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 31.0992 LAYER M4 ;
  END BIAS_ADJ[2]
  PIN BIAS_ADJ[1] 
    ANTENNAPARTIALMETALAREA 0.054 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
  END BIAS_ADJ[1]
  PIN BIAS_ADJ[0] 
    ANTENNAPARTIALMETALAREA 0.0595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
  END BIAS_ADJ[0]
  PIN BIAS_DBP[13] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M3 ;
  END BIAS_DBP[13]
  PIN BIAS_DBP[12] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0655 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3322 LAYER M2 ;
  END BIAS_DBP[12]
  PIN BIAS_DBP[11] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.342 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9488 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.82 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 47.696 LAYER M6 ;
  END BIAS_DBP[11]
  PIN BIAS_DBP[10] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.4495 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0218 LAYER M3 ;
  END BIAS_DBP[10]
  PIN BIAS_DBP[9] 
    ANTENNAPARTIALMETALAREA 0.099 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4356 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.266 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2144 LAYER M3 ;
  END BIAS_DBP[9]
  PIN BIAS_DBP[8] 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DBP[8]
  PIN BIAS_DBP[7] 
    ANTENNAPARTIALMETALAREA 0.378 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7072 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.1328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.422 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.5008 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.218 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0032 LAYER M6 ;
  END BIAS_DBP[7]
  PIN BIAS_DBP[6] 
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.438 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9712 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.782 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.2848 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.758 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 42.9792 LAYER M6 ;
  END BIAS_DBP[6]
  PIN BIAS_DBP[5] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.104 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5016 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.358 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 50.1072 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 264.497 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1169.31 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA6 ;
  END BIAS_DBP[5]
  PIN BIAS_DBP[4] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.438 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.5712 LAYER M4 ;
  END BIAS_DBP[4]
  PIN BIAS_DBP[3] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.698 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1152 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 3.982 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.5648 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.736 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 47.3264 LAYER M6 ;
  END BIAS_DBP[3]
  PIN BIAS_DBP[2] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.218 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.718 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.0032 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.338 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.5312 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 503.071 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2220.43 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_DBP[2]
  PIN BIAS_DBP[1] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.558 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.702 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5328 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.754 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 51.8496 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 0.246 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1264 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M7 ; 
    ANTENNAMAXAREACAR 63.934 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 284.926 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA7 ;
  END BIAS_DBP[1]
  PIN BIAS_DBP[0] 
    ANTENNAPARTIALMETALAREA 0.0225 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.882 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7248 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.062 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 44.3168 LAYER M6 ;
  END BIAS_DBP[0]
  PIN BIAS_DBN[13] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6528 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.666 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3744 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 8.158 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 35.9392 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 185.343 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 817.864 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.2987 LAYER VIA6 ;
  END BIAS_DBN[13]
  PIN BIAS_DBN[12] 
    ANTENNAPARTIALMETALAREA 2.2205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.8142 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.338 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3312 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.586 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4224 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.702 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3328 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 122.255 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 540.277 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_DBN[12]
  PIN BIAS_DBN[11] 
    ANTENNAPARTIALMETALAREA 0.061 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2684 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.548 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.542 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 33.2288 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 185.783 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 820.563 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_DBN[11]
  PIN BIAS_DBN[10] 
    ANTENNAPARTIALMETALAREA 3.1315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.566 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.118 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 22.5632 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 112.666 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 498.323 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.0101 LAYER VIA6 ;
  END BIAS_DBN[10]
  PIN BIAS_DBN[9] 
    ANTENNAPARTIALMETALAREA 0.258 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1792 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0608 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 2.182 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.6448 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.058 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 26.6992 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 178.983 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 790.643 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA6 ;
  END BIAS_DBN[9]
  PIN BIAS_DBN[8] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.082 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 2.246 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9264 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.818 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.4432 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 196.183 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 867.057 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA6 ;
  END BIAS_DBN[8]
  PIN BIAS_DBN[7] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.668 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.5167 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 69.9233 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.5 LAYER VIA3 ;
  END BIAS_DBN[7]
  PIN BIAS_DBN[6] 
    ANTENNAPARTIALMETALAREA 2.6295 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5698 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7024 LAYER M3 ;
  END BIAS_DBN[6]
  PIN BIAS_DBN[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.796 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.2784 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.522 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3408 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.976 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.5824 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 0.382 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M7 ; 
    ANTENNAMAXAREACAR 73.6254 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 328.835 LAYER M7 ;
    ANTENNAMAXCUTCAR 3.23625 LAYER VIA7 ;
  END BIAS_DBN[5]
  PIN BIAS_DBN[4] 
    ANTENNAPARTIALMETALAREA 0.0625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.275 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.098 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8752 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 1.286 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7024 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.976 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 26.3824 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 0.784 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5376 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER M7 ; 
    ANTENNAMAXAREACAR 56.1311 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 250.764 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.56695 LAYER VIA7 ;
  END BIAS_DBN[4]
  PIN BIAS_DBN[3] 
    ANTENNAPARTIALMETALAREA 0.057 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2508 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.52 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.0224 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 62.1097 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.577201 LAYER VIA3 ;
  END BIAS_DBN[3]
  PIN BIAS_DBN[2] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
  END BIAS_DBN[2]
  PIN BIAS_DBN[1] 
    ANTENNAPARTIALMETALAREA 0.022 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.854 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2456 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.072 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3608 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.062 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7168 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 2.696 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 11.9504 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 215.151 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 949.411 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA6 ;
  END BIAS_DBN[1]
  PIN BIAS_DBN[0] 
    ANTENNAPARTIALMETALAREA 0.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.818 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0432 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.582 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.2048 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.886 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 8.3424 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.898 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5952 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 328.391 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1449.18 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.589 LAYER VIA6 ;
  END BIAS_DBN[0]
  PIN BIAS_DBPC[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.219 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0076 LAYER M2 ;
  END BIAS_DBPC[13]
  PIN BIAS_DBPC[12] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_DBPC[12]
  PIN BIAS_DBPC[11] 
    ANTENNAPARTIALMETALAREA 0.126 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5544 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.338 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5312 LAYER M3 ;
  END BIAS_DBPC[11]
  PIN BIAS_DBPC[10] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.1355 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6402 LAYER M2 ;
  END BIAS_DBPC[10]
  PIN BIAS_DBPC[9] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.692 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1328 LAYER M3 ;
  END BIAS_DBPC[9]
  PIN BIAS_DBPC[8] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.6885 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0734 LAYER M3 ;
  END BIAS_DBPC[8]
  PIN BIAS_DBPC[7] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
  END BIAS_DBPC[7]
  PIN BIAS_DBPC[6] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 11.288 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 49.7552 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 3.462 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 15.2768 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 90.591 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 400.003 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.94175 LAYER VIA7 ;
  END BIAS_DBPC[6]
  PIN BIAS_DBPC[5] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 5.382 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.7248 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 3.74 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 16.544 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 97.7886 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 432.332 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.443 LAYER VIA6 ;
  END BIAS_DBPC[5]
  PIN BIAS_DBPC[4] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5648 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 10.334 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 45.6016 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 0.226 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0384 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M7 ; 
    ANTENNAMAXAREACAR 107.796 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 481.217 LAYER M7 ;
    ANTENNAMAXCUTCAR 3.55987 LAYER VIA7 ;
  END BIAS_DBPC[4]
  PIN BIAS_DBPC[3] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.136 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.1632 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.378 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.7072 LAYER M6 ;
  END BIAS_DBPC[3]
  PIN BIAS_DBPC[2] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.258 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2232 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.058 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.742 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.1088 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 457.768 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2020.98 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.23625 LAYER VIA6 ;
  END BIAS_DBPC[2]
  PIN BIAS_DBPC[1] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.342 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.898 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9952 LAYER M4 ;
  END BIAS_DBPC[1]
  PIN BIAS_DBPC[0] 
    ANTENNAPARTIALMETALAREA 0.5805 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5982 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.606 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1104 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.542 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.2288 LAYER M4 ;
  END BIAS_DBPC[0]
  PIN BIAS_DBNC[13] 
    ANTENNAPARTIALMETALAREA 0.055 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 2.938 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9712 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.102 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.0928 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 203.104 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 897.276 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_DBNC[13]
  PIN BIAS_DBNC[12] 
    ANTENNAPARTIALMETALAREA 0.4485 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9734 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.466 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4944 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 6.758 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 29.7792 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M6 ; 
    ANTENNAMAXAREACAR 150.168 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 664.99 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.1544 LAYER VIA6 ;
  END BIAS_DBNC[12]
  PIN BIAS_DBNC[11] 
    ANTENNAPARTIALMETALAREA 0.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 3.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 9.942 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 43.7888 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 234.601 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1036.06 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_DBNC[11]
  PIN BIAS_DBNC[10] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 3.598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8752 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5984 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.968 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.176 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4624 LAYER M6 ;
  END BIAS_DBNC[10]
  PIN BIAS_DBNC[9] 
    ANTENNAPARTIALMETALAREA 0.053 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.678 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4272 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 3.678 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.2272 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.106 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.968 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 4.918 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.6832 LAYER M6 ;
  END BIAS_DBNC[9]
  PIN BIAS_DBNC[8] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1232 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.162 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7568 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 10.158 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 44.7392 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 1.766 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 7.8144 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M7 ; 
    ANTENNAMAXAREACAR 56.0342 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 250.37 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.66667 LAYER VIA7 ;
  END BIAS_DBNC[8]
  PIN BIAS_DBNC[7] 
    ANTENNAPARTIALMETALAREA 0.051 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2244 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.746 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7704 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.052 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 2.498 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 11.0352 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 65.7675 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 292.463 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.33333 LAYER VIA6 ;
  END BIAS_DBNC[7]
  PIN BIAS_DBNC[6] 
    ANTENNAPARTIALMETALAREA 0.0565 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2486 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4752 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.622 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1808 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M5 ; 
    ANTENNAMAXAREACAR 157.534 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 696.237 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA5 ;
  END BIAS_DBNC[6]
  PIN BIAS_DBNC[5] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.686 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2992 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 5.302 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.3728 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.078 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 22.3872 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 455.485 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2009.4 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.91262 LAYER VIA6 ;
  END BIAS_DBNC[5]
  PIN BIAS_DBNC[4] 
    ANTENNAPARTIALMETALAREA 0.1445 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6358 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.138 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8512 LAYER M4 ;
  END BIAS_DBNC[4]
  PIN BIAS_DBNC[3] 
    ANTENNAPARTIALMETALAREA 0.076 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.498 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8352 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 82.4621 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 365.18 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA4 ;
  END BIAS_DBNC[3]
  PIN BIAS_DBNC[2] 
    ANTENNAPARTIALMETALAREA 1.7525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.755 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.306 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M3 ;
  END BIAS_DBNC[2]
  PIN BIAS_DBNC[1] 
    ANTENNAPARTIALMETALAREA 0.088 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.286 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M3 ;
  END BIAS_DBNC[1]
  PIN BIAS_DBNC[0] 
    ANTENNAPARTIALMETALAREA 0.0195 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.032 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.098 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8752 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.626 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1984 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 5.5 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 24.288 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M6 ; 
    ANTENNAMAXAREACAR 257.505 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1139.94 LAYER M6 ;
    ANTENNAMAXCUTCAR 2.589 LAYER VIA6 ;
  END BIAS_DBNC[0]
  PIN BIAS_TC_POT[5] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.2475 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.133 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.998 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4352 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 20.7675 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 92.9967 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA4 ;
  END BIAS_TC_POT[5]
  PIN BIAS_TC_POT[4] 
    ANTENNAPARTIALMETALAREA 0.575 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.53 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.722 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2208 LAYER M3 ;
  END BIAS_TC_POT[4]
  PIN BIAS_TC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.8045 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.346 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.5675 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.45 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.662 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3568 LAYER M4 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 52.2675 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 233.063 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA4 ;
  END BIAS_TC_POT[3]
  PIN BIAS_TC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.486 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1384 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.9008 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 48.85 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.222 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.8208 LAYER M4 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 47.9342 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 212.53 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA4 ;
  END BIAS_TC_POT[2]
  PIN BIAS_TC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.211 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9284 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0775 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.385 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.586 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6224 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 55.2654 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 244.874 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.809061 LAYER VIA4 ;
  END BIAS_TC_POT[1]
  PIN BIAS_TC_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.062 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.678 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.0032 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 62.6084 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.485437 LAYER VIA3 ;
  END BIAS_TC_POT[0]
  PIN BIAS_LC_POT[5] 
    ANTENNAPARTIALMETALAREA 0.111 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4884 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.006 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.0167 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 106.59 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3872 LAYER M4 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 25.3167 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 113.043 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M5 ;
    ANTENNAGATEAREA 0.06 LAYER M5 ; 
    ANTENNAMAXAREACAR 26.65 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 119.643 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.598 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0752 LAYER M6 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 53.2833 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 237.563 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_LC_POT[5]
  PIN BIAS_LC_POT[4] 
    ANTENNAPARTIALMETALAREA 0.224 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9856 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.502 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2528 LAYER M3 ;
  END BIAS_LC_POT[4]
  PIN BIAS_LC_POT[3] 
    ANTENNAPARTIALMETALAREA 0.8115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6146 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.314 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.15 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 32.3767 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.118 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5632 LAYER M4 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 9.11667 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 41.7633 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAMAXCUTCAR 1.16667 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 0.106 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5104 LAYER M5 ;
    ANTENNAGATEAREA 0.06 LAYER M5 ; 
    ANTENNAMAXAREACAR 10.8833 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 50.27 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 2.158 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 9.5392 LAYER M6 ;
    ANTENNAGATEAREA 0.06 LAYER M6 ; 
    ANTENNAMAXAREACAR 46.85 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 209.257 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.5 LAYER VIA6 ;
  END BIAS_LC_POT[3]
  PIN BIAS_LC_POT[2] 
    ANTENNAPARTIALMETALAREA 0.192 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1856 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.464 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.3296 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 LAYER M4 ; 
    ANTENNAMAXAREACAR 65.95 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 292.563 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA4 ;
  END BIAS_LC_POT[2]
  PIN BIAS_LC_POT[1] 
    ANTENNAPARTIALMETALAREA 0.047 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.6325 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.827 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.408 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 56.248 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 249.699 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.61812 LAYER VIA4 ;
  END BIAS_LC_POT[1]
  PIN BIAS_LC_POT[0] 
    ANTENNAPARTIALMETALAREA 0.306 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.442 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9888 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 12.2876 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 55.534 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.809061 LAYER VIA4 ;
  END BIAS_LC_POT[0]
  PIN BIAS_TIA_G_POT[15] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2078 LAYER M2 ;
  END BIAS_TIA_G_POT[15]
  PIN BIAS_TIA_G_POT[14] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.529 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3716 LAYER M2 ;
  END BIAS_TIA_G_POT[14]
  PIN BIAS_TIA_G_POT[13] 
    ANTENNAPARTIALMETALAREA 0.6525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.871 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.618 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7632 LAYER M3 ;
  END BIAS_TIA_G_POT[13]
  PIN BIAS_TIA_G_POT[12] 
    ANTENNAPARTIALMETALAREA 0.397 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7468 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.446 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.2064 LAYER M3 ;
  END BIAS_TIA_G_POT[12]
  PIN BIAS_TIA_G_POT[11] 
    ANTENNAPARTIALMETALAREA 0.611 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6884 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.162 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1568 LAYER M3 ;
  END BIAS_TIA_G_POT[11]
  PIN BIAS_TIA_G_POT[10] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.289 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2716 LAYER M2 ;
  END BIAS_TIA_G_POT[10]
  PIN BIAS_TIA_G_POT[9] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1525 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.115 LAYER M2 ;
  END BIAS_TIA_G_POT[9]
  PIN BIAS_TIA_G_POT[8] 
    ANTENNAPARTIALMETALAREA 0.176 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M3 ;
  END BIAS_TIA_G_POT[8]
  PIN BIAS_TIA_G_POT[7] 
    ANTENNAPARTIALMETALAREA 1.7125 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.535 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.426 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9184 LAYER M3 ;
  END BIAS_TIA_G_POT[7]
  PIN BIAS_TIA_G_POT[6] 
    ANTENNAPARTIALMETALAREA 0.107 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4708 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.958 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2592 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 15.102 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 66.4928 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0893 LAYER M5 ; 
    ANTENNAMAXAREACAR 187.791 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 824.591 LAYER M5 ;
    ANTENNAMAXCUTCAR 0.895857 LAYER VIA5 ;
  END BIAS_TIA_G_POT[6]
  PIN BIAS_TIA_G_POT[5] 
    ANTENNAPARTIALMETALAREA 0.0695 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3058 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.462 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4768 LAYER M5 ;
  END BIAS_TIA_G_POT[5]
  PIN BIAS_TIA_G_POT[4] 
    ANTENNAPARTIALMETALAREA 0.335 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.474 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.702 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1328 LAYER M3 ;
  END BIAS_TIA_G_POT[4]
  PIN BIAS_TIA_G_POT[3] 
    ANTENNADIFFAREA 1.458 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.5455 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4442 LAYER M2 ;
  END BIAS_TIA_G_POT[3]
  PIN BIAS_TIA_G_POT[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.816 LAYER M2 ;
  END BIAS_TIA_G_POT[2]
  PIN BIAS_TIA_G_POT[1] 
    ANTENNAPARTIALMETALAREA 0.6345 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7918 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.926 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5184 LAYER M3 ;
  END BIAS_TIA_G_POT[1]
  PIN BIAS_TIA_G_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.922 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1008 LAYER M2 ;
  END BIAS_TIA_G_POT[0]
  PIN BIAS_REV_POT[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.154 LAYER M2 ;
  END BIAS_REV_POT[13]
  PIN BIAS_REV_POT[12] 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.658 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9392 LAYER M4 ;
  END BIAS_REV_POT[12]
  PIN BIAS_REV_POT[11] 
    ANTENNAPARTIALMETALAREA 0.182 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8008 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.746 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3264 LAYER M3 ;
  END BIAS_REV_POT[11]
  PIN BIAS_REV_POT[10] 
    ANTENNAPARTIALMETALAREA 0.0235 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1034 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
  END BIAS_REV_POT[10]
  PIN BIAS_REV_POT[9] 
    ANTENNAPARTIALMETALAREA 0.062 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.738 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.0912 LAYER M4 ;
  END BIAS_REV_POT[9]
  PIN BIAS_REV_POT[8] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.3745 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0918 LAYER M2 ;
  END BIAS_REV_POT[8]
  PIN BIAS_REV_POT[7] 
    ANTENNAPARTIALMETALAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.378 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7072 LAYER M3 ;
  END BIAS_REV_POT[7]
  PIN BIAS_REV_POT[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.038 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M2 ;
  END BIAS_REV_POT[6]
  PIN BIAS_REV_POT[5] 
    ANTENNAPARTIALMETALAREA 0.072 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3168 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.862 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8368 LAYER M3 ;
  END BIAS_REV_POT[5]
  PIN BIAS_REV_POT[4] 
    ANTENNAPARTIALMETALAREA 0.1375 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.605 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9568 LAYER M3 ;
  END BIAS_REV_POT[4]
  PIN BIAS_REV_POT[3] 
    ANTENNAPARTIALMETALAREA 0.025 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.11 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.762 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3968 LAYER M3 ;
  END BIAS_REV_POT[3]
  PIN BIAS_REV_POT[2] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.4625 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.123 LAYER M2 ;
  END BIAS_REV_POT[2]
  PIN BIAS_REV_POT[1] 
    ANTENNAPARTIALMETALAREA 0.058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2552 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.402 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M3 ;
  END BIAS_REV_POT[1]
  PIN BIAS_REV_POT[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4158 LAYER M2 ;
  END BIAS_REV_POT[0]
  PIN BIAS_TC_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.191 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8404 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.7295 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2538 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.948 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6592 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 31.4538 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 139.72 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA4 ;
  END BIAS_TC_DSADC[5]
  PIN BIAS_TC_DSADC[4] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.368 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0632 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.186 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.838 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.3312 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 18.042 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 79.4288 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNADIFFAREA 1.696 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.138 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6512 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNADIFFAREA 1.696 LAYER M7 ; 
    ANTENNAPARTIALMETALAREA 10.732 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 47.3968 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M7 ; 
    ANTENNAMAXAREACAR 210.41 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 931.489 LAYER M7 ;
    ANTENNAMAXCUTCAR 1.45631 LAYER VIA7 ;
  END BIAS_TC_DSADC[4]
  PIN BIAS_TC_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.1645 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7238 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.362 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6368 LAYER M3 ;
  END BIAS_TC_DSADC[3]
  PIN BIAS_TC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0693 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.30231 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 27.1371 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.486 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1824 LAYER M4 ;
    ANTENNAGATEAREA 0.0693 LAYER M4 ; 
    ANTENNAMAXAREACAR 13.3153 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 58.6291 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.721501 LAYER VIA4 ;
  END BIAS_TC_DSADC[2]
  PIN BIAS_TC_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.1775 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.781 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.966 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2944 LAYER M3 ;
  END BIAS_TC_DSADC[1]
  PIN BIAS_TC_DSADC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.708 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1592 LAYER M2 ;
  END BIAS_TC_DSADC[0]
  PIN BIAS_LC_DSADC[5] 
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1935 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8954 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.788 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5552 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M4 ; 
    ANTENNAMAXAREACAR 40.4167 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 180.777 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA4 ;
  END BIAS_LC_DSADC[5]
  PIN BIAS_LC_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.797 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.21 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M3 ; 
    ANTENNAMAXAREACAR 81.1088 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 358.489 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA3 ;
  END BIAS_LC_DSADC[4]
  PIN BIAS_LC_DSADC[3] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.8941 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.971 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.542 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.102 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.318 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.2432 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 52.4098 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 232.146 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA5 ;
  END BIAS_LC_DSADC[3]
  PIN BIAS_LC_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.087 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3828 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.0828 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.678 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0272 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 3.076 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.6224 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 62.3451 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 270.476 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.2945 LAYER VIA5 ;
  END BIAS_LC_DSADC[2]
  PIN BIAS_LC_DSADC[1] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.9845 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4198 LAYER M2 ;
  END BIAS_LC_DSADC[1]
  PIN BIAS_LC_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.699 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0756 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.022 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5408 LAYER M3 ;
  END BIAS_LC_DSADC[0]
  PIN BIAS_RIN_DSADC[5] 
    ANTENNAPARTIALMETALAREA 0.5325 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.343 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.078 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.1872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 82.6828 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 365.023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER VIA3 ;
  END BIAS_RIN_DSADC[5]
  PIN BIAS_RIN_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7172 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.322 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4608 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.942 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5888 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 50.7087 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 220.667 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA5 ;
  END BIAS_RIN_DSADC[4]
  PIN BIAS_RIN_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.091 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.182 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 0.962 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2768 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M5 ; 
    ANTENNAMAXAREACAR 57.1748 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 253.987 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.13269 LAYER VIA5 ;
  END BIAS_RIN_DSADC[3]
  PIN BIAS_RIN_DSADC[2] 
    ANTENNAPARTIALMETALAREA 0.612 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6928 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0208 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6288 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 LAYER M4 ; 
    ANTENNAMAXAREACAR 19.9903 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 90.3754 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.809061 LAYER VIA4 ;
  END BIAS_RIN_DSADC[2]
  PIN BIAS_RIN_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.2505 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1022 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.848 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 LAYER M3 ; 
    ANTENNAMAXAREACAR 99.1877 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 439.068 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.970874 LAYER VIA3 ;
  END BIAS_RIN_DSADC[1]
  PIN BIAS_RIN_DSADC[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.43 LAYER M2 ;
  END BIAS_RIN_DSADC[0]
  PIN BIAS_RFB_DSADC[5] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.955 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.29 LAYER M2 ;
  END BIAS_RFB_DSADC[5]
  PIN BIAS_RFB_DSADC[4] 
    ANTENNAPARTIALMETALAREA 0.457 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0108 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.298 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3552 LAYER M3 ;
  END BIAS_RFB_DSADC[4]
  PIN BIAS_RFB_DSADC[3] 
    ANTENNAPARTIALMETALAREA 0.8105 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8928 LAYER M3 ;
  END BIAS_RFB_DSADC[3]
  PIN BIAS_RFB_DSADC[2] 
    ANTENNAPARTIALMETALAREA 1.965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.646 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.682 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4448 LAYER M3 ;
  END BIAS_RFB_DSADC[2]
  PIN BIAS_RFB_DSADC[1] 
    ANTENNAPARTIALMETALAREA 0.711 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1284 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.658 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9392 LAYER M3 ;
  END BIAS_RFB_DSADC[1]
  PIN BIAS_RFB_DSADC[0] 
    ANTENNAPARTIALMETALAREA 0.655 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.002 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4528 LAYER M3 ;
  END BIAS_RFB_DSADC[0]
  PIN BIAS_DSADC_VCM[13] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 3.677 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.1788 LAYER M2 ;
  END BIAS_DSADC_VCM[13]
  PIN BIAS_DSADC_VCM[12] 
    ANTENNAPARTIALMETALAREA 0.0555 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.918 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0832 LAYER M4 ;
  END BIAS_DSADC_VCM[12]
  PIN BIAS_DSADC_VCM[11] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6752 LAYER M4 ;
  END BIAS_DSADC_VCM[11]
  PIN BIAS_DSADC_VCM[10] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.102 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4928 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.038 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6112 LAYER M4 ;
  END BIAS_DSADC_VCM[10]
  PIN BIAS_DSADC_VCM[9] 
    ANTENNAPARTIALMETALAREA 3.581 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8004 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNADIFFAREA 1.696 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.278 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6672 LAYER M4 ;
  END BIAS_DSADC_VCM[9]
  PIN BIAS_DSADC_VCM[8] 
    ANTENNAPARTIALMETALAREA 0.0535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.142 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6688 LAYER M3 ;
  END BIAS_DSADC_VCM[8]
  PIN BIAS_DSADC_VCM[7] 
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.692 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.282 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2848 LAYER M3 ;
  END BIAS_DSADC_VCM[7]
  PIN BIAS_DSADC_VCM[6] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.0585 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3014 LAYER M2 ;
  END BIAS_DSADC_VCM[6]
  PIN BIAS_DSADC_VCM[5] 
    ANTENNAPARTIALMETALAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2596 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.662 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9568 LAYER M3 ;
  END BIAS_DSADC_VCM[5]
  PIN BIAS_DSADC_VCM[4] 
    ANTENNAPARTIALMETALAREA 0.0205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.042 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6288 LAYER M3 ;
  END BIAS_DSADC_VCM[4]
  PIN BIAS_DSADC_VCM[3] 
    ANTENNAPARTIALMETALAREA 0.189 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8316 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.742 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3088 LAYER M3 ;
  END BIAS_DSADC_VCM[3]
  PIN BIAS_DSADC_VCM[2] 
    ANTENNAPARTIALMETALAREA 0.0965 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.458 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.822 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6608 LAYER M3 ;
  END BIAS_DSADC_VCM[2]
  PIN BIAS_DSADC_VCM[1] 
    ANTENNAPARTIALMETALAREA 0.031 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.738 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2912 LAYER M3 ;
  END BIAS_DSADC_VCM[1]
  PIN BIAS_DSADC_VCM[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.3075 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.397 LAYER M2 ;
  END BIAS_DSADC_VCM[0]
  PIN dsadc_conv_done 
    ANTENNAPARTIALMETALAREA 0.106 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4664 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 10.938 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.1712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M3 ; 
    ANTENNAMAXAREACAR 469.945 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 2064.83 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.63265 LAYER VIA3 ;
  END dsadc_conv_done
  PIN dsadc_en 
    ANTENNAPARTIALMETALAREA 1.262 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5528 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1968 LAYER M3 ;
  END dsadc_en
  PIN dsadc_clk 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.224 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3224 LAYER M3 ;
  END dsadc_clk
  PIN dsadc_switch[2] 
    ANTENNAPARTIALMETALAREA 0.5495 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.842 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.5488 LAYER M3 ;
  END dsadc_switch[2]
  PIN dsadc_switch[1] 
    ANTENNAPARTIALMETALAREA 0.271 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.399 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.1996 LAYER M3 ;
  END dsadc_switch[1]
  PIN dsadc_switch[0] 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 1.1595 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1018 LAYER M2 ;
  END dsadc_switch[0]
  PIN dac_en_pot 
    ANTENNADIFFAREA 1.696 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.346 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5664 LAYER M2 ;
  END dac_en_pot
  PIN adc_ext_in 
    ANTENNAPARTIALMETALAREA 0.107 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4708 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.482 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.5648 LAYER M3 ;
  END adc_ext_in
  PIN atp_en 
    ANTENNAPARTIALMETALAREA 0.3205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4102 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.422 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 1.058 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6992 LAYER M5 ;
  END atp_en
  PIN atp_sel 
    ANTENNAPARTIALMETALAREA 0.375 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.65 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.522 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.3408 LAYER M3 ;
  END atp_sel
  PIN adc_sel 
    ANTENNAPARTIALMETALAREA 0.2095 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9218 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.686 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0624 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.202 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9328 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNADIFFAREA 1.696 LAYER M5 ; 
    ANTENNAPARTIALMETALAREA 2.978 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.1472 LAYER M5 ;
  END adc_sel
  PIN saradc_clk 
    ANTENNAPARTIALMETALAREA 1.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNADIFFAREA 1.696 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 70.462 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.0362 LAYER M3 ;
  END saradc_clk
  PIN saradc_rdy 
    ANTENNAPARTIALMETALAREA 0.7715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3946 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8304 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.402 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8128 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.738 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 60.4912 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M5 ; 
    ANTENNAMAXAREACAR 503.801 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2220.54 LAYER M5 ;
    ANTENNAMAXCUTCAR 1.72911 LAYER VIA5 ;
  END saradc_rdy
  PIN saradc_rst 
    ANTENNADIFFAREA 1.692 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 0.2915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER M2 ;
  END saradc_rst
  PIN saradc_data[9] 
    ANTENNAPARTIALMETALAREA 0.1825 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.803 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.052 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2728 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.566 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5344 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.698 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 60.3152 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M5 ; 
    ANTENNAMAXAREACAR 455.187 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 1994.83 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.30548 LAYER VIA5 ;
  END saradc_data[9]
  PIN saradc_data[8] 
    ANTENNAPARTIALMETALAREA 0.047 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2068 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1735 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8074 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.926 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1184 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.038 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 57.4112 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0271 LAYER M5 ; 
    ANTENNAMAXAREACAR 547.223 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2414.44 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.58303 LAYER VIA5 ;
  END saradc_data[8]
  PIN saradc_data[7] 
    ANTENNAPARTIALMETALAREA 0.4315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.306 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3904 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.338 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.5312 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.146 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6864 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6 ; 
    ANTENNAMAXAREACAR 481.412 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2127.08 LAYER M6 ;
    ANTENNAMAXCUTCAR 3.67347 LAYER VIA6 ;
  END saradc_data[7]
  PIN saradc_data[6] 
    ANTENNAPARTIALMETALAREA 0.7115 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1306 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.1444 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3344 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.396 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 5.698 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 25.1152 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.166 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7744 LAYER M6 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA6 ;
    ANTENNAPARTIALMETALAREA 2.234 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9616 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0347 LAYER M7 ; 
    ANTENNAMAXAREACAR 154.092 LAYER M7 ;
    ANTENNAMAXSIDEAREACAR 686.726 LAYER M7 ;
    ANTENNAMAXCUTCAR 2.88184 LAYER VIA7 ;
  END saradc_data[6]
  PIN saradc_data[5] 
    ANTENNAPARTIALMETALAREA 0.8915 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9226 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.538 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3024 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 6.576 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 29.0224 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA5 ;
    ANTENNAPARTIALMETALAREA 0.372 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M6 ; 
    ANTENNAMAXAREACAR 202.271 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 899.576 LAYER M6 ;
    ANTENNAMAXCUTCAR 4.08163 LAYER VIA6 ;
  END saradc_data[5]
  PIN saradc_data[4] 
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.7135 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1834 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.826 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6784 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 9.296 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.9904 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 560.067 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2468.56 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[4]
  PIN saradc_data[3] 
    ANTENNAPARTIALMETALAREA 0.8715 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8346 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.278 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6672 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.526 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3584 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.938 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 61.3712 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 678.745 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2988.33 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[3]
  PIN saradc_data[2] 
    ANTENNAPARTIALMETALAREA 1.0315 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5386 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6704 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.302 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.638 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 60.0512 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 637.673 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2811.32 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.85714 LAYER VIA5 ;
  END saradc_data[2]
  PIN saradc_data[1] 
    ANTENNAPARTIALMETALAREA 0.427 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8788 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.01 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 0.5535 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4794 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.206 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9504 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.98 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 61.6 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 644.965 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2835.31 LAYER M5 ;
    ANTENNAMAXCUTCAR 3.26531 LAYER VIA5 ;
  END saradc_data[1]
  PIN saradc_data[0] 
    ANTENNAPARTIALMETALAREA 0.771 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA2 ;
    ANTENNAPARTIALMETALAREA 1.0935 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8554 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 0.104 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5016 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.02 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 13.616 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 59.9984 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 LAYER M5 ; 
    ANTENNAMAXAREACAR 647.512 LAYER M5 ;
    ANTENNAMAXSIDEAREACAR 2850.4 LAYER M5 ;
    ANTENNAMAXCUTCAR 2.85714 LAYER VIA5 ;
  END saradc_data[0]
END MCU

END LIBRARY
